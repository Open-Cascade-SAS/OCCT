-- Created on: 1995-06-20
-- Created by: Stagiaire Alain JOURDAIN <ajo@phobox>
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class IncrementalMesh from BRepMesh

inherits DiscretRoot from BRepMesh

    ---Purpose: Builds the mesh of a shape with respect of their
    --          correctly triangulated parts
    --

uses
    Box from Bnd,
    Shape from TopoDS,
    Face  from TopoDS,
    Edge  from TopoDS,
    MapOfShape  from TopTools,
    IndexedDataMapOfShapeListOfShape from TopTools,
    DataMapOfShapeReal from TopTools,
    FastDiscret  from BRepMesh,
    Status       from BRepMesh,
    PDiscretRoot from BRepMesh

is
    Create
        returns IncrementalMesh from BRepMesh;
    ---C++: alias "Standard_EXPORT virtual ~BRepMesh_IncrementalMesh();"

    Create (S       : Shape   from TopoDS;
            D       : Real    from Standard;
            Relatif : Boolean from Standard = Standard_False;
            Ang     : Real    from Standard = 0.5)
        returns IncrementalMesh from BRepMesh;
    ---Purpose: If the  boolean    <Relatif>   is  True,    the
    --          deflection used   for the polygonalisation   of
    --          each edge will be <D> * Size of Edge.
    --          the deflection used for the faces will be the maximum
    --          deflection of their edges.

    SetRelative (     me : mutable;
                 theFlag : Boolean from Standard);

    Relative (me)
        returns Boolean from Standard;

    Init (me : mutable)
        is redefined protected;

    Perform (me : mutable)
        is redefined;

    Update (me : mutable;
             S : Shape from TopoDS)
        is static;
    ---Purpose: Builds the incremental mesh of the shape

    IsModified (me)
        returns Boolean from Standard
        is static;

    Update (me : mutable;
            E  : Edge from TopoDS)
        is static private;
    ---Purpose: Locate a correct discretisation if it exists
    --          Set no one otherwise

    Update (me : mutable;
            F  : Face from TopoDS)
        is static private;
    ---Purpose: If the face is  not correctly triangulated, or
    --          if  one  of its edges  is  to be discretisated
    --          correctly, the triangulation  of this face  is
    --          built.

    GetStatusFlags (me)
        returns Integer from Standard
        is static;

    SetParallel (           me : mutable;
                 theInParallel : Boolean from Standard);
    ---Purpose:
    -- Request algorithm to launch in multiple threads to improve performance.

    IsParallel (me)
        returns Boolean from Standard;
    ---Purpose:
    -- Returns the multi-threading usage flag.

    --
    --  Plugin interface
    --
    Discret (myclass;
             theShape      : Shape from TopoDS;
             theDeflection : Real from Standard;
             theAngle      : Real from Standard;
             theAlgo       : out PDiscretRoot from BRepMesh)
        returns Integer from Standard;
    ---Purpose:
    -- Plugin interface for the Mesh Factories.

    IsParallelDefault (myclass)
        returns Boolean from Standard;
    ---Purpose:
    -- Returns multi-threading usage flag set by default in
    -- Discret() static method (thus applied only to Mesh Factories).

    SetParallelDefault (myclass;
                        theInParallel : Boolean from Standard);
    ---Purpose:
    -- Setup multi-threading usage flag set by default in
    -- Discret() static method (thus applied only to Mesh Factories).

fields
    myRelative   : Boolean     from Standard is protected;
    myInParallel : Boolean     from Standard is protected;
    myMap        : MapOfShape  from TopTools is protected;
    myMesh       : FastDiscret from BRepMesh is protected;
    myModified   : Boolean     from Standard is protected;
    mymapedge    : DataMapOfShapeReal from TopTools is protected;
    myancestors  : IndexedDataMapOfShapeListOfShape from TopTools is protected;
    mydtotale    : Real from Standard is protected;
    myBox        : Box  from Bnd is protected;
    myStatus     : Integer from Standard is protected;

end IncrementalMesh;
