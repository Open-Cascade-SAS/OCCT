-- File:	RWStepDimTol_RWConcentricityTolerance.cdl
-- Created:	Wed Jun  4 13:34:34 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWConcentricityTolerance from RWStepDimTol

    ---Purpose: Read & Write tool for ConcentricityTolerance

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ConcentricityTolerance from StepDimTol

is
    Create returns RWConcentricityTolerance from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ConcentricityTolerance from StepDimTol);
	---Purpose: Reads ConcentricityTolerance

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ConcentricityTolerance from StepDimTol);
	---Purpose: Writes ConcentricityTolerance

    Share (me; ent : ConcentricityTolerance from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWConcentricityTolerance;
