-- Created on: 1999-09-08
-- Created by: Andrey BETENEV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class MeasureRepresentationItem from StepRepr 
    inherits RepresentationItem from StepRepr 

	---Purpose: Implements a measure_representation_item entity
	--          which is used for storing validation properties
	--          (e.g. area) for shapes

uses
    HAsciiString       from TCollection,
    Unit               from StepBasic,
    MeasureWithUnit    from StepBasic,
    MeasureValueMember from StepBasic
    
is
    Create returns mutable MeasureRepresentationItem;
        ---Purpose: Creates empty object
    
    Init (me : mutable;
	  aName : mutable HAsciiString from TCollection;
	  aValueComponent : MeasureValueMember from StepBasic;
	  aUnitComponent : Unit from StepBasic);
        ---Purpose: Init all fields

    SetMeasure (me: mutable; Measure: MeasureWithUnit from StepBasic);
    Measure (me) returns MeasureWithUnit from StepBasic;
    
fields
    myMeasure: MeasureWithUnit from StepBasic;

end MeasureRepresentationItem;

