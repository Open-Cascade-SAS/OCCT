-- File:	StepFEA_NodeRepresentation.cdl
-- Created:	Thu Dec 12 17:51:06 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class NodeRepresentation from StepFEA
inherits Representation from StepRepr

    ---Purpose: Representation of STEP entity NodeRepresentation

uses
    HAsciiString from TCollection,
    HArray1OfRepresentationItem from StepRepr,
    RepresentationContext from StepRepr,
    FeaModel from StepFEA

is
    Create returns NodeRepresentation from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aRepresentation_Name: HAsciiString from TCollection;
                       aRepresentation_Items: HArray1OfRepresentationItem from StepRepr;
                       aRepresentation_ContextOfItems: RepresentationContext from StepRepr;
                       aModelRef: FeaModel from StepFEA);
	---Purpose: Initialize all fields (own and inherited)

    ModelRef (me) returns FeaModel from StepFEA;
	---Purpose: Returns field ModelRef
    SetModelRef (me: mutable; ModelRef: FeaModel from StepFEA);
	---Purpose: Set field ModelRef

fields
    theModelRef: FeaModel from StepFEA;

end NodeRepresentation;
