-- Created on: 2002-10-29
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package BinLDrivers

uses
    Standard,
    TDF,
    TCollection,
    TColStd,
    CDM,
    PCDM,
    Storage,
    BinObjMgt,
    BinMDF

is

    class DocumentStorageDriver;
    class DocumentRetrievalDriver;

    class    DocumentSection;
    imported VectorOfDocumentSection;

    Factory (theGUID : GUID from Standard) returns Transient from Standard;

    AttributeDrivers (MsgDrv : MessageDriver from CDM)
        returns ADriverTable from BinMDF;
        ---Purpose: Creates a table of the supported drivers' types

    StorageVersion returns AsciiString from TCollection;
        ---Purpose: returns last storage version
    
end BinLDrivers;
