-- Created on: 1993-06-22
-- Created by: Jean Louis FRENKEL
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



-- Modified:	Jeudi 26 Janvier 1995
-- by:		CAL
--		The old name of this was Marker.

deferred class VectorialMarker from Graphic2d inherits Line from Graphic2d

	---Version:

	---Purpose: Groups all the primitives which behaves like
	--	    geometrical marker.
	--	    for example : EllipsMarker, CircleMarker ...
	--	    A marker is a primitive which retains its original
	--	    on-screen size no matter how the view is zoomed.
	--	    For example, markers are used as symbols of dimension.
	--	    Every marker takes a reference point as an argument in
	--	    its constructor. CircleMarker and EllipsMarker take
	--	    another point as the center and PolylineMarker takes the
	--	    first point of its list as its origin.
	--	    The coordinates of the centre or origin point are offsets
	--	    with respect to the reference point.

	---Keywords: Primitive, VectorialMarker
	---Warning:
	---References:

uses
	GraphicObject	from Graphic2d,
	Length		from Quantity

is
	-------------------------
	-- Category: Constructors
	-------------------------

	Initialize (aGraphicObject: GraphicObject from Graphic2d;
		aXPosition, aYPosition: Length from Quantity);
	---Level: Public
	---Purpose: Creates a marker at <aXPosition>, <aYPosition>
	---Category: Constructors

	---------------------------------------------------
	-- Category: Methods to modify the class definition
	---------------------------------------------------

	SetPosition (me: mutable;
		aXPosition, aYPosition: Length from Quantity)
	is static;
	---Level: Public
	---Purpose: Modifies the marker position.
	--  Warning: If the associated GraphicObject is transformed
	--	    the position will be transformed.
	---Category: Methods to modify the class definition

	----------------------------
	-- Category: Inquire methods
	----------------------------

	XPosition (me) returns Length from Quantity
	is static;
	---Level: Public
	---Purpose: Returns the x position of the marker
	--  Warning: If the associated GraphicObject is transformed
	--	    the returned position is the transformed position.
	---Category: Inquire methods

	YPosition (me) returns Length from Quantity is static;
	---Level: Public
	---Purpose: Returns the y position of the marker
	--  Warning: If the associated GraphicObject is transformed
	--	    the returned position is the transformed position.
	---Category: Inquire methods

fields
	myXPosition:	ShortReal from Standard is protected;
	myYPosition:	ShortReal from Standard is protected;

end VectorialMarker from Graphic2d;
