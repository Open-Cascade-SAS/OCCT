-- File:	RWStepDimTol_RWDatumTarget.cdl
-- Created:	Wed Jun  4 13:34:35 2003 
-- Author:	Galina KULIKOVA
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWDatumTarget from RWStepDimTol

    ---Purpose: Read & Write tool for DatumTarget

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    DatumTarget from StepDimTol

is
    Create returns RWDatumTarget from RWStepDimTol;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : DatumTarget from StepDimTol);
	---Purpose: Reads DatumTarget

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: DatumTarget from StepDimTol);
	---Purpose: Writes DatumTarget

    Share (me; ent : DatumTarget from StepDimTol;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWDatumTarget;
