-- Created on: 1995-01-05
-- Created by: Frederic MAUPAS
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class GeometricTool from StepToTopoDS

  ---Purpose: This class contains some algorithmic services 
  --          specific to the mapping STEP to CAS.CADE              

uses

    Tool         from StepToTopoDS,
    SurfaceCurve from StepGeom,
    Surface      from StepGeom,
    Pcurve       from StepGeom,
    EdgeLoop     from StepShape,    
    Edge         from StepShape,    
    Curve        from Geom2d,
    Line         from Geom2d,
    Curve        from Geom,
    Surface      from Geom,
    Pnt2d        from gp,
    Pnt          from gp,
    Face         from TopoDS,
    Wire         from TopoDS,
    Edge         from TopoDS,
    Vertex       from TopoDS
    
is

    PCurve(myclass;
 	      SC : SurfaceCurve from StepGeom;
    	      S  : Surface      from StepGeom;
	      PC : out Pcurve   from StepGeom;
	      last : Integer = 0)
    	returns Integer;

    IsSeamCurve(myclass;
    	    	SC : SurfaceCurve from StepGeom;
    	      	S  : Surface      from StepGeom;
		E  : Edge         from StepShape;
    	    	EL : EdgeLoop     from StepShape)
    	returns Boolean;

		
    IsLikeSeam(myclass;
    	       SC : SurfaceCurve from StepGeom;
       	       S  : Surface      from StepGeom;
	       E  : Edge         from StepShape;
    	       EL : EdgeLoop     from StepShape)
    	returns Boolean;


    UpdateParam3d(myclass; C  : Curve from Geom;
    	    	  w1, w2 : in out Real from Standard;
		  preci  : Real)
    	returns Boolean;
			 
end GeometricTool from StepToTopoDS;
