-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( Kiran )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TransformationMatrix from IGESGeom  inherits TransfEntity

        ---Purpose: defines IGESTransformationMatrix, Type <124> Form <0>
        --          in package IGESGeom
        --          The transformation matrix entity transforms three-row column
        --          vectors by means of matrix multiplication and then a vector
        --          addition. This entity can be considered as an "operator"
        --          entity in that it starts with the input vector, operates on
        --          it as described above, and produces the output vector.

uses

        HArray2OfReal from TColStd,
	IGESEntity    from IGESData,
        GTrsf         from gp

raises DimensionMismatch, OutOfRange

is

        Create returns mutable TransformationMatrix;

        -- Specific Methods pertaining to the class

        Init (me      : mutable;
              aMatrix : HArray2OfReal)
        raises DimensionMismatch;
        ---Purpose : This method is used to set the fields of the class
        --           TransformationMatrix
        --       - aMatrix : 3 x 4 array containing elements of the
        --                   transformation matrix
        -- raises exception if aMatrix is not 3 x 4 array

    	SetFormNumber (me : mutable; form : Integer) raises OutOfRange;
	---Purpose : Changes FormNumber (indicates the Type of Transf :
	--           Transformation 0-1 or Coordinate System 10-11-12)
	--           Error if not in ranges [0-1] or [10-12]

    	Data (me; I, J : Integer) returns Real  raises OutOfRange;
	---Purpose : returns individual Data
	-- Errro if I not in [1-3] or J not in [1-4]


        Value (me) returns GTrsf;
        ---Purpose : returns the transformation matrix
        -- 4th row elements of GTrsf will always be 0, 0, 0, 1 (not defined)

fields

--
-- Class    : IGESGeom_TransformationMatrix
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class TransformationMatrix.
--
-- Reminder : A TransformationMatrix instance is defined by :
--            the coefficients of a 3 X 4 matrix

        theData : HArray2OfReal;

end TransformationMatrix;
