-- File:	RWStepBasic_RWContract.cdl
-- Created:	Fri Nov 26 16:26:37 1999 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class RWContract from RWStepBasic

    ---Purpose: Read & Write tool for Contract

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    Contract from StepBasic

is
    Create returns RWContract from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : Contract from StepBasic);
	---Purpose: Reads Contract

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: Contract from StepBasic);
	---Purpose: Writes Contract

    Share (me; ent : Contract from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWContract;
