-- Created on: 1992-05-15
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class InteriorPoint from IntSurf

	---Purpose: Definition of a point solution of the
	--          intersection between an implicit an a
	--          parametrised surface. These points are
	--          passing points on the intersection lines,
	--          or starting points for the closed lines
	--          on the parametrised surface.


uses Pnt   from gp,
     Vec   from gp,
     Vec2d from gp

is

    Create
    
    	returns InteriorPoint from IntSurf;


    Create(P: Pnt from gp; U,V: Real from Standard;
           Direc: Vec from gp; Direc2d: Vec2d from gp)
	   
	returns InteriorPoint from IntSurf;


    SetValue(me: in out; P: Pnt from gp; U,V: Real from Standard;
           Direc: Vec from gp; Direc2d: Vec2d from gp)
	   
	is static;


    Value(me)
    
	---Purpose: Returns the 3d coordinates of the interior point.

    	returns Pnt from gp
    	---C++: return const&
	---C++: inline

	is static;


    Parameters(me; U,V: out Real from Standard)
    
	---Purpose: Returns the parameters of the interior point on the
	--          parametric surface.
    
	---C++: inline

    	is static;


    UParameter(me)
    
	---Purpose: Returns the first parameter of the interior point on the
	--          parametric surface.

    	returns Real from Standard
	---C++: inline
    
    	is static;


    VParameter(me)
    
	---Purpose: Returns the second parameter of the interior point on the
	--          parametric surface.
    
    	returns Real from Standard
	---C++: inline
    
    	is static;


    Direction(me)

        ---Purpose: Returns the tangent at the intersection in 3d space
        --          associated to the interior point.
    
    	returns Vec from gp
    	---C++: return const&
	---C++: inline
	
	is static;


    Direction2d(me)

        ---Purpose: Returns the tangent at the intersection in the parametric
        --          space of the parametric surface.
    
    	returns Vec2d from gp
    	---C++: return const&
	---C++: inline
	
	is static;

fields

    point   : Pnt   from gp;
    paramu  : Real  from Standard;
    paramv  : Real  from Standard;
    direc   : Vec   from gp;
    direc2d : Vec2d from gp;

end InteriorPoint;
