-- Created on: 1997-01-08
-- Created by: VAUTHIER Jean-Claude
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



package QADNaming 

	---Purpose: 

	--           FOR OLD TOPOLOGY ONLY!
uses 
    Draw,
    TCollection, 
    TColStd,
    TDF,
    TNaming,
    TopoDS,
    TopTools
is
         
    class DataMapOfShapeOfName instantiates
    	DataMap from TCollection(Shape          from TopoDS,
	    	    	    	 AsciiString    from TCollection,
                                 ShapeMapHasher from TopTools);  				  			       								   
    CurrentShape (ShapeEntry      : CString  from Standard; 
    	    	  Data            : Data     from TDF)
    returns Shape from TopoDS;		  

    GetShape (ShapeEntry  :        CString     from Standard; 
    	      Data        :        Data        from TDF;
    	      Shapes      : in out ListOfShape from TopTools);
    

    GetEntry (Shape      : in     Shape   from TopoDS; 
              Data       : in     Data    from TDF; 
              Status     : in out Integer from Standard)
    	---Purpose: Status = 0  Not  found, 
    	--          Status = 1  One  shape,
    	--          Status = 2  More than one shape. 
    returns AsciiString from TCollection;
    
    Entry (theArguments : Address from Standard;
    	   theLabel : in out Label from TDF) returns Boolean from Standard;
    --- Purpose: returns label by first two arguments (df and entry string)

    AllCommands        (DI : in out Interpretor from Draw);
    
    BasicCommands      (DI : in out Interpretor from Draw);
    ---Purpose: commands relatives to NamedShape

    BuilderCommands    (DI : in out Interpretor from Draw);
    ---Purpose: loading NamedShape to the Data Framework

    IteratorsCommands  (DI : in out Interpretor from Draw);
    ---Purpose: loading NamedShape to the Data Framework

    ToolsCommands      (DI : in out Interpretor from Draw);
    
    SelectionCommands  (DI : in out Interpretor from Draw);
    ---Purpose: commands relatives to Naming 

end QADNaming;




