-- Created on: 1997-08-07
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Session from CDF inherits Transient from Standard


uses
    Directory from CDF,
    ExtendedString from TCollection,
    Application from CDF, 
    MetaDataDriver from CDF, 
    Writer from PCDM
raises

    NoSuchObject from Standard,MultiplyDefined from Standard

is
    Create  returns mutable Session from CDF
    raises MultiplyDefined from Standard;

    Exists(myclass)
--- Purpose: returns true if a session has been created.
    returns Boolean from Standard;
    
    CurrentSession(myclass) returns mutable Session from CDF;
    ---Purpose: returns the only one instance of Session 
    --          that has been created.

    
    Directory(me) returns mutable Directory from CDF;
    ---Purpose: returns the directory of the session;
    ---Level: Public 

    
---Category: current application management
    HasCurrentApplication(me) returns Boolean from Standard;
    
    CurrentApplication(me) returns mutable Application from CDF
    raises NoSuchObject from Standard;
    
    SetCurrentApplication(me: mutable; anApplication: Application from CDF);
    
    UnsetCurrentApplication(me: mutable);


---Category: database related methods

    MetaDataDriver(me) returns MetaDataDriver from CDF
    raises NoSuchObject from Standard;
    
    
    LoadDriver(me: mutable);

fields

    myDirectory            : Directory from CDF;
    myCurrentApplication   : Application from CDF;
    myHasCurrentApplication: Boolean from Standard;
    myMetaDataDriver       : MetaDataDriver from CDF;
friends
    class Application from CDF
end Session from CDF;
