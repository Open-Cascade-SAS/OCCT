-- Created on: 1994-04-18
-- Created by: Modelistation
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Marker2D from Draw inherits Drawable2D from Draw

	---Purpose: 

uses
    Pnt2d from gp,
    Color from Draw,
    MarkerShape from Draw,
    Display from Draw

is
    Create(P : Pnt2d from gp; T : MarkerShape from Draw; C : Color from Draw; 
    	Size : Integer = 5) returns mutable Marker2D from Draw;
	
    Create(P : Pnt2d from gp; T : MarkerShape from Draw; C : Color from Draw; 
    	RSize : Real) returns mutable Marker2D from Draw;
    
    ChangePos(me : mutable) returns Pnt2d from gp;
    ---C++: return &
    ---Purpose: myPos field

    DrawOn(me; dis : in out Display from Draw);

    PickReject(me; X,Y,Prec : Real) returns Boolean
	---Purpose: Returs always false
    is redefined;
    

fields
    myPos : Pnt2d from gp;
    myCol : Color from Draw;
    myTyp : MarkerShape from Draw;
    mySiz : Integer;

end Marker2D;
