-- File:	RWStepBasic_RWExternalSource.cdl
-- Created:	Wed May 10 15:09:06 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.1
-- Copyright:	Matra Datavision 2000

class RWExternalSource from RWStepBasic

    ---Purpose: Read & Write tool for ExternalSource

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    ExternalSource from StepBasic

is
    Create returns RWExternalSource from RWStepBasic;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : ExternalSource from StepBasic);
	---Purpose: Reads ExternalSource

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: ExternalSource from StepBasic);
	---Purpose: Writes ExternalSource

    Share (me; ent : ExternalSource from StepBasic;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWExternalSource;
