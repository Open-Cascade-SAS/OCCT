-- Created on: 1999-10-01
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 1999-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ImportShape from QANewBRepNaming inherits TopNaming from QANewBRepNaming

    ---Purpose: This class provides a topological naming 
    --          of a Shape

uses 
 
    Shape     from TopoDS,
    Label     from TDF,
    LabelMap  from TDF,
    TagSource from TDF

is 
 
    Create returns ImportShape from QANewBRepNaming;    

    Create (ResultLabel : Label from TDF) 
    returns ImportShape from QANewBRepNaming;  

    Init (me : in out; ResultLabel : Label from TDF);
    

    Load (me; S : Shape from TopoDS);
    ---Purpose: Use this method for a topological naming of a Shape

    LoadPrime (me; S : Shape from TopoDS);

    LoadFirstLevel (me; S : Shape from TopoDS; Tagger : TagSource from TDF);

    LoadNextLevels (me; S : Shape from TopoDS; Tagger : TagSource from TDF);

    LoadC0Edges(me; S : Shape from TopoDS; 
    	     	       Tagger : TagSource from TDF);
    ---Purpose: Method for internal use. It is used by Load().
    --          It loads the edges which couldn't be uniquely identified as 
    --          an intersection of two faces.


    LoadC0Vertices (me; S : Shape from TopoDS; Tagger : TagSource from TDF);

    NamedFaces (me; theNamedFaces : in out LabelMap from TDF)
    returns Integer from Standard;

    NamedEdges (me; theNamedEdges : in out LabelMap from TDF)
    returns Integer from Standard;

    NamedVertices (me; theNamedVertices : in out LabelMap from TDF)
    returns Integer from Standard;

end ImportShape;	       
