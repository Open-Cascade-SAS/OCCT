-- Created on: 1997-02-24
-- Created by: Olga PILLOT
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Revol from LocOpe 

	---Purpose: Defines a prism (using Prism from BRepSweep)
	--          with modifications provided for the Prism feature.

 
uses DataMapOfShapeListOfShape from TopTools,
     ListOfShape               from TopTools,
     Ax1                       from gp,     
     Shape from TopoDS,
     SequenceOfCurve from TColGeom, 
     Curve            from  Geom, 
     Vec              from  gp
     

raises NoSuchObject from Standard,
       NotDone      from StdFail

is

 
    Create 
     
    	returns  Revol  from  LocOpe;


    Create (Base     : Shape   from  TopoDS;
    	    Axis     : Ax1     from  gp;
    	    Angle    : Real    from  Standard;
    	    angledec : Real    from  Standard)
	    
	returns Revol from LocOpe;     

    Create (Base   : Shape from TopoDS;
    	    Axis     : Ax1     from  gp;
    	    Angle    : Real    from  Standard)

	returns Revol from LocOpe;     


    Perform(me:  in  out;  Base     : Shape   from  TopoDS; 
	        	   Axis     : Ax1     from  gp;
    	    	    	   Angle    : Real    from  Standard;
    	                   angledec : Real    from  Standard)
			    
	is  static;


    Perform(me:  in  out;  Base     :  Shape  from  TopoDS; 
	        	   Axis     : Ax1     from  gp;
    	    	    	   Angle    : Real    from  Standard) 
			    
	is  static;


    FirstShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    LastShape(me)
    
    	returns Shape from TopoDS
	---C++: return const &
	is static;


    Shape(me)
    
    	returns Shape from TopoDS 
	raises  NotDone  from  StdFail
	---C++: return const &
	is static;


    Shapes(me; S: Shape from TopoDS)
    
    	returns ListOfShape from TopTools
	---C++: return const &
    	raises NoSuchObject from Standard
	       -- The exception is raised if S is not a subshape of the profile
	is static;


    Curves(me;  SCurves:  in  out  SequenceOfCurve  from  TColGeom)
    
	is static;
 

    BarycCurve(me) 
     
    	returns  Curve  from  Geom 
	is  static;
  
    IntPerf(me:  in  out) 
     
    	is  static  private;
 

fields

    myBase       : Shape             from  TopoDS;
    myAxis       : Ax1               from  gp; 
    myAngle      : Real              from  Standard; 
    myAngTra     : Real              from  Standard;
    myIsTrans    : Boolean           from  Standard;
    myDone       : Boolean           from  Standard; 
    myRes        : Shape             from  TopoDS;
    myFirstShape : Shape             from  TopoDS;
    myLastShape  : Shape             from  TopoDS;
    myMap        : DataMapOfShapeListOfShape    from TopTools;
     
end Prism;     
