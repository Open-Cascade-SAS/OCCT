-- File:	RWStepFEA_RWFeaAreaDensity.cdl
-- Created:	Thu Dec 12 17:51:05 2002 
-- Author:	data exchange team
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2
-- Copyright:	Open CASCADE 2002

class RWFeaAreaDensity from RWStepFEA

    ---Purpose: Read & Write tool for FeaAreaDensity

uses
    Check from Interface,
    StepWriter from StepData,
    StepReaderData from StepData,
    EntityIterator from Interface,
    FeaAreaDensity from StepFEA

is
    Create returns RWFeaAreaDensity from RWStepFEA;
	---Purpose: Empty constructor

    ReadStep (me; data: StepReaderData from StepData; num: Integer;
                  ach : in out Check from Interface;
                  ent : FeaAreaDensity from StepFEA);
	---Purpose: Reads FeaAreaDensity

    WriteStep (me; SW: in out StepWriter from StepData;
                   ent: FeaAreaDensity from StepFEA);
	---Purpose: Writes FeaAreaDensity

    Share (me; ent : FeaAreaDensity from StepFEA;
               iter: in out EntityIterator from Interface);
	---Purpose: Fills data for graph (shared items)

end RWFeaAreaDensity;
