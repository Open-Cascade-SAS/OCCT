-- Created on: 2003-02-04
-- Created by: data exchange team
-- Copyright (c) 2003-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class ElementGeometricRelationship from StepFEA
inherits TShared from MMgt

    ---Purpose: Representation of STEP entity ElementGeometricRelationship

uses
    ElementOrElementGroup from StepFEA,
    AnalysisItemWithinRepresentation from StepElement,
    ElementAspect from StepElement

is
    Create returns ElementGeometricRelationship from StepFEA;
	---Purpose: Empty constructor

    Init (me: mutable; aElementRef: ElementOrElementGroup from StepFEA;
                       aItem: AnalysisItemWithinRepresentation from StepElement;
                       aAspect: ElementAspect from StepElement);
	---Purpose: Initialize all fields (own and inherited)

    ElementRef (me) returns ElementOrElementGroup from StepFEA;
	---Purpose: Returns field ElementRef
    SetElementRef (me: mutable; ElementRef: ElementOrElementGroup from StepFEA);
	---Purpose: Set field ElementRef

    Item (me) returns AnalysisItemWithinRepresentation from StepElement;
	---Purpose: Returns field Item
    SetItem (me: mutable; Item: AnalysisItemWithinRepresentation from StepElement);
	---Purpose: Set field Item

    Aspect (me) returns ElementAspect from StepElement;
	---Purpose: Returns field Aspect
    SetAspect (me: mutable; Aspect: ElementAspect from StepElement);
	---Purpose: Set field Aspect

fields
    theElementRef: ElementOrElementGroup from StepFEA;
    theItem: AnalysisItemWithinRepresentation from StepElement;
    theAspect: ElementAspect from StepElement;

end ElementGeometricRelationship;
