-- Created on: 1997-10-01
-- Created by: Christian CAILLET
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SelectFaces  from IGESSelect  inherits SelectExplore

    ---Purpose : This selection returns the faces contained in an IGES Entity
    --           or itself if it is a Face
    --           Face means :
    --           - Face (510) of a ManifoldSolidBrep
    --           - TrimmedSurface (144)
    --           - BoundedSurface (143)
    --           - Plane with a Bounding Curve (108, form not 0)
    --           - Also, any Surface which is not in a TrimmedSurface, a
    --             BoundedSurface, or a Face (FREE Surface)
    --           -> i.e. a Face for which Natural Bounds will be considered

uses AsciiString from TCollection, Transient, EntityIterator, Graph

is


    Create returns mutable  SelectFaces;


    Explore (me; level : Integer; ent : Transient; G : Graph;
    	     explored : in out EntityIterator)
    	returns Boolean;
    ---Purpose : Explores an entity, to take its faces
    --           Works recursively


    ExploreLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns a text defining the criterium : "Faces"

end SelectFaces;
