-- Created on: 2002-12-12
-- Created by: data exchange team
-- Copyright (c) 2002-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.2

class SymmetricTensor22d from StepFEA
inherits SelectType from StepData

    ---Purpose: Representation of STEP SELECT type SymmetricTensor22d

uses
    HArray1OfReal from TColStd

is
    Create returns SymmetricTensor22d from StepFEA;
	---Purpose: Empty constructor

    CaseNum (me; ent: Transient) returns Integer;
	---Purpose: Recognizes a kind of SymmetricTensor22d select type
	--          1 -> HArray1OfReal from TColStd
	--          0 else

    AnisotropicSymmetricTensor22d (me) returns HArray1OfReal from TColStd;
	---Purpose: Returns Value as AnisotropicSymmetricTensor22d (or Null if another type)

end SymmetricTensor22d;
