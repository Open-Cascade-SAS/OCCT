-- Created on: 1991-03-06
-- Created by: Denis Pascal
-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

generic class VertexIterator from GraphTools (Graph  as any;
		    		               Vertex as any)
				  
--template class VertexIterator from GraphTools (Graph  as any,
--                                                 Vertex as any)
				  
    ---Purpose: Template class which  defines Signature of an iterator
    --          to visit each adjacent vertex  of a  given one  in the
    --          underlying graph.


raises NoMoreObject from Standard,
       NoSuchObject from Standard

is

    Create (G : Graph; V : Vertex) returns VertexIterator;

    More (me) returns Boolean;
	---Purpose: Returns TRUE if there are other vertices.
       ---Level: Public

    Next(me : in out)
    	--- Purpose : Set the iterator to the next Vertex.
       ---Level: Public
    raises NoMoreObject from Standard;

    Value(me) returns Vertex
	--- Purpose: Returns the vertex value for the current position
	--           of the iterator.
       ---Level: Public
    raises NoSuchObject from Standard;

end VertexIterator;



















