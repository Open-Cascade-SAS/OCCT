-- Created on: 1995-08-25
-- Created by: Remi LEQUETTE
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class HSurface from GeomAdaptor inherits GHSurface from GeomAdaptor

    	---Purpose: An interface between the services provided by any
    	-- surface from the package Geom and those required
    	-- of the surface by algorithms which use it.

uses
    Surface from Geom,
    Surface from GeomAdaptor

raises
    ConstructionError from Standard

is

    Create returns mutable HSurface from GeomAdaptor;
    	---C++: inline
    
    Create( AS : Surface from GeomAdaptor) returns mutable HSurface from GeomAdaptor;
    	---C++: inline

    Create( S : Surface from Geom) returns mutable HSurface from GeomAdaptor;
    	---C++: inline
    
    Create( S : Surface from Geom; UFirst,ULast,VFirst,VLast : Real; 
    	    TolU  :  Real  =  0.0; 
            TolV  :  Real  =  0.0) 
    returns  mutable HSurface from GeomAdaptor
    raises ConstructionError from Standard;
    	---Purpose: ConstructionError is raised if UFirst>ULast or VFirst>VLast
    	---C++: inline

end HSurface;
