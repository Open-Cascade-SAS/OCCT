-- Created on: 1994-08-03
-- Created by: Christophe MARION
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Algo from HLRBRep inherits InternalAlgo from HLRBRep

    	---Purpose: A framework to compute a shape as seen in a projection plane. This is done by
    	-- calculating the visible and the hidden parts of the shape.
    	-- HLRBRep_Algo works with three types of entity:
    	-- -   shapes to be visualized
    	-- -   edges in these shapes (these edges are
    	-- the basic entities which will be visualized or hidden), and
    	-- -   faces in these shapes which hide the edges.
    	--   HLRBRep_Algo is based on the principle of comparing each edge of the shape to be
    	-- visualized with each of its faces, and calculating the visible and the hidden parts of each edge.
    	-- For a given projection, HLRBRep_Algo calculates a set of lines characteristic of the
    	-- object being represented. It is also used in conjunction with the
    	-- HLRBRep_HLRToShape extraction utilities, which reconstruct a new, simplified shape
    	-- from a selection of calculation results. This new shape is made up of edges, which
    	-- represent the shape visualized in the projection.
    	-- HLRBRep_Algo takes the shape itself into account whereas HLRBRep_PolyAlgo
    	-- works with a polyhedral simplification of the shape. When you use HLRBRep_Algo, you
    	-- obtain an exact result, whereas, when you use HLRBRep_PolyAlgo, you reduce
    	-- computation time but obtain polygonal segments. In the case of complicated
    	-- shapes, HLRBRep_Algo may be time-consuming.
    	-- An HLRBRep_Algo object provides a framework for:
    	-- -   defining the point of view
    	-- -   identifying the shape or shapes to be visualized
    	-- -   calculating the outlines
    	-- -   calculating the visible and hidden lines of the shape.
    	--   Warning
    	-- -   Superimposed lines are not eliminated by this algorithm.
    	-- -   There must be no unfinished objects inside the shape you wish to visualize.
    	-- -   Points are not treated.
    	-- -   Note that this is not the sort of algorithm used in generating shading, which
    	--   calculates the visible and hidden parts of each face in a shape to be visualized by
    	--   comparing each face in the shape with every other face in the same shape.
        
uses
    TShared from MMgt,
    Shape   from TopoDS

is
    Create returns mutable Algo from HLRBRep;
    	---Purpose: Constructs an empty framework for the
    	-- calculation of visible and hidden lines of a shape in a projection.
    	-- Use the function:
    	-- -   Projector to define the point of view
    	-- -   Add to select the shape or shapes to be visualized
    	-- -   Update to compute the outlines of the shape, and
    	-- -   Hide to compute the visible and hidden lines of the shape.
    
    Create(A : Algo from HLRBRep) returns mutable Algo from HLRBRep;

    Add(me : mutable; S     : Shape   from TopoDS;
    	    	      SData : TShared from MMgt;
                      nbIso : Integer from Standard = 0)
	---Purpose: add the Shape <S>.
    is static;
    
    Add(me : mutable; S     : Shape   from TopoDS;
                      nbIso : Integer from Standard = 0)
	---Purpose:  Adds the shape S to this framework, and
    	-- specifies the number of isoparameters nbiso desired in visualizing S.
    	-- You may add as many shapes as you wish. Use the function Add once for each shape.
    is static;
    
    Index(me : mutable; S : Shape from TopoDS)
    returns Integer from Standard
	---Purpose: return  the index  of  the  Shape <S>  and
	--          return 0 if the Shape <S> is not found.
    is static;

    OutLinedShapeNullify(me : mutable)
	---Purpose: nullify all the results of OutLiner from HLRTopoBRep.
    is static;
    
end Algo;
