-- File:	MeshAlgo_Triangle.cdl
-- Created:	Tue May 11 16:43:27 1993
-- Author:	Didier PIFFAULT
--		<dpf@nonox>
---Copyright:	 Matra Datavision 1993

-- signature
deferred class Triangle from MeshAlgo

	---Purpose: Describes the   data structure of  a  Triangle for
	--          Deleaunay triangulation.


uses    Boolean from Standard,
    	Integer from Standard,
    	ListOfInteger from TColStd,
	DegreeOfFreedom from MeshDS


is      Initialize     (e1, e2, e3 : Integer from Standard;
	    	    	o1, o2, o3 : Boolean from Standard;
                        canMove : DegreeOfFreedom from MeshDS);
    	
	
	Edges          (me;
	    	    	e1, e2, e3 : out Integer from Standard;
	    	    	o1, o2, o3 : out Boolean from Standard);


    	Movability     (me)
    	    returns DegreeOfFreedom from MeshDS;


	SetMovability  (me      : in out;
    	    	    	   canMove : DegreeOfFreedom from MeshDS);


---Purpose: For maping the Triangles.
--          Same Triangle -> Same HashCode
--          Different Triangles -> Not IsEqual but can have same HashCode 

    	HashCode      (me;
    	    	       Upper : Integer from Standard)
	---C++: function call
    	        returns Integer from Standard;


    	IsEqual       (me; Other : Triangle from MeshAlgo)
	---C++: alias operator ==
	    returns Boolean from Standard;

end Triangle;
