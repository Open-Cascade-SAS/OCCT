-- Created on: 1993-11-16
-- Created by: Laurent BOURESCHE
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class FaceInterference from ChFiDS 

	---Purpose: interference face/fillet

uses Curve from Geom2d,
     Orientation from TopAbs

is
    Create returns FaceInterference from ChFiDS;
    
    SetInterference(me             : in out; 
    	    	    LineIndex      : Integer from Standard;
		    Trans          : Orientation from TopAbs; 
    	    	    PCurv1 ,PCurv2 : Curve from Geom2d )is static;
    ---C++: inline
    	    	
    SetTransition(me : in out; Trans : Orientation from TopAbs) is static;
    
    SetFirstParameter(me : in out; U1 : Real)    is static;
    ---C++: inline
    	    	
    SetLastParameter(me : in out; U1 : Real)     is static;
    ---C++: inline
    	    	
    SetParameter(me      : in out; 
    	    	 U1      : Real from Standard;
                 IsFirst : Boolean from Standard)
    is static;
  
    LineIndex(me) returns Integer from Standard;
    ---C++: inline
    	    	
    SetLineIndex(me : in out; I : Integer from Standard);
    ---C++: inline
    	    	
    Transition(me) returns Orientation from TopAbs is static;
    ---C++: inline

    PCurveOnFace(me) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return const &

    PCurveOnSurf(me) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return const &

    ChangePCurveOnFace(me : in out) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return &

    ChangePCurveOnSurf(me : in out) returns Curve from Geom2d is static;
    ---C++: inline
    ---C++: return &

    FirstParameter(me) returns Real from Standard is static ;
    ---C++: inline

    LastParameter(me) returns Real from Standard is static;
    ---C++: inline

    Parameter(me; IsFirst : Boolean from Standard) 
    returns Real from Standard is static;

fields

firstParam     : Real        from Standard;
lastParam      : Real        from Standard;
pCurveOnFace   : Curve       from Geom2d;
pCurveOnSurf   : Curve       from Geom2d; 
lineindex      : Integer     from Standard;
LineTransition : Orientation from TopAbs;
end FaceInterference;
