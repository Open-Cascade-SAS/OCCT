-- Created on: 2000-05-24
-- Created by: Edward AGAPOV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class DocumentRetrievalDriver from XCAFDrivers 
inherits DocumentRetrievalDriver from MDocStd

	---Purpose: retrieval driver of a XS document

uses
    ARDriverTable from MDF,
    MessageDriver from CDM

is
    Create returns DocumentRetrievalDriver from XCAFDrivers;    

    AttributeDrivers(me : mutable; theMessageDriver : MessageDriver from CDM)
    returns ARDriverTable from MDF
    is redefined;

end DocumentRetrievalDriver;

