-- File:	MDataStd_RealArrayRetrievalDriver.cdl
-- Created:	Tue Jun 15 16:56:00 1999
-- Author:	Sergey RUIN
---Copyright:	 Matra Datavision 1999


class RealArrayRetrievalDriver from MDataStd inherits ARDriver from MDF

	---Purpose: 

uses RRelocationTable from MDF,
     Attribute        from TDF,
     Attribute        from PDF, 
     MessageDriver    from CDM
is

    Create(theMessageDriver : MessageDriver from CDM)  -- Version 0
    returns mutable RealArrayRetrievalDriver from MDataStd;


    VersionNumber(me) returns Integer from Standard;
	---Purpose: Returns the version number from which the driver
	--          is available: 0.

    SourceType(me) returns Type from Standard;
	---Purpose: Returns the type: RealArray from PDataStd.

    NewEmpty (me) returns mutable Attribute from TDF;


    Paste(me;
    	  Source     :         Attribute from PDF;
    	  Target     : mutable Attribute from TDF;
    	  RelocTable : RRelocationTable from MDF);


end RealArrayRetrievalDriver;

