-- Copyright (c) 1991-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Dir2d    from gp   inherits Storable

        ---Purpose: Describes a unit vector in the plane (2D space). This unit
        -- vector is also called "Direction".
        -- See Also
        -- gce_MakeDir2d which provides functions for more
        -- complex unit vector constructions
        -- Geom2d_Direction which provides additional functions
        -- for constructing unit vectors and works, in particular, with
        -- the parametric equations of unit vectors

uses  Ax2d   from gp,
      Trsf2d from gp,
      Vec2d  from gp,
      XY     from gp

raises ConstructionError from Standard,
       DomainError       from Standard,
       OutOfRange        from Standard


is


 
  Create  returns Dir2d;
        --- Purpose : Creates a direction corresponding to X axis.
    	---C++:inline
   
  Create (V : Vec2d)  returns Dir2d
        --- Purpose : Normalizes the vector V and creates a Direction. Raises ConstructionError if V.Magnitude() <= Resolution from gp.
    	---C++:inline
     raises ConstructionError;
   
  Create (Coord : XY)   returns Dir2d
        --- Purpose : Creates a Direction from a doublet of coordinates. Raises ConstructionError if Coord.Modulus() <= Resolution from gp.
    	---C++:inline
     raises ConstructionError;

  Create ( Xv, Yv : Real)  returns Dir2d
        --- Purpose : Creates a Direction with its 2 cartesian coordinates. Raises ConstructionError if Sqrt(Xv*Xv + Yv*Yv) <= Resolution from gp.
    	---C++:inline
     raises ConstructionError;
       
  SetCoord (me: in out; Index : Integer; Xi : Real)
    	---C++:inline  
        --- Purpose :
    	--      For this unit vector, assigns:
    	-- the value Xi to:
    	--   -   the X coordinate if Index is 1, or
    	--   -   the Y coordinate if Index is 2, and then normalizes it.
    	-- Warning
    	-- Remember that all the coordinates of a unit vector are
    	-- implicitly modified when any single one is changed directly.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is not 1 or 2.
    	-- Standard_ConstructionError if either of the following
    	-- is less than or equal to gp::Resolution():
    	-- -   Sqrt(Xv*Xv + Yv*Yv), or
    	-- -   the modulus of the number pair formed by the new
    	--   value Xi and the other coordinate of this vector that
    	--   was not directly modified.   
        --  Raises OutOfRange if Index != {1, 2}.
     raises OutOfRange,
            ConstructionError
     is static;

  SetCoord (me : in out; Xv, Yv : Real)  raises ConstructionError  is static;
    	---C++:inline  
        --- Purpose :
    	--      For this unit vector, assigns:
    	-- -   the values Xv and Yv to its two coordinates, 
    	-- Warning
    	-- Remember that all the coordinates of a unit vector are
    	-- implicitly modified when any single one is changed directly.
    	-- Exceptions
    	-- Standard_OutOfRange if Index is not 1 or 2.
    	-- Standard_ConstructionError if either of the following
    	-- is less than or equal to gp::Resolution():
    	-- -   Sqrt(Xv*Xv + Yv*Yv), or
    	-- -   the modulus of the number pair formed by the new
    	--   value Xi and the other coordinate of this vector that
    	--   was not directly modified.   
    	--  Raises OutOfRange if Index != {1, 2}.   

  SetX (me: in out; X : Real)            raises ConstructionError  is static;
    	---C++:inline  
    	---Purpose:
    	-- Assigns the given value to the X coordinate of this unit   vector,
    	--   and then normalizes it.
    	-- Warning
    	-- Remember that all the coordinates of a unit vector are
    	-- implicitly modified when any single one is changed directly.
    	-- Exceptions
    	-- Standard_ConstructionError if either of the following
    	-- is less than or equal to gp::Resolution():
    	-- -   the modulus of Coord, or
    	-- -   the modulus of the number pair formed from the new
    	--   X or Y coordinate and the other coordinate of this
    	--   vector that was not directly modified.

  SetY (me: in out; Y : Real)            raises ConstructionError  is static;
    	---C++:inline  
    	---Purpose:
    	-- Assigns  the given value to the Y coordinate of this unit   vector,
    	--   and then normalizes it.
    	-- Warning
    	-- Remember that all the coordinates of a unit vector are
    	-- implicitly modified when any single one is changed directly.
    	-- Exceptions
    	-- Standard_ConstructionError if either of the following
    	-- is less than or equal to gp::Resolution():
    	-- -   the modulus of Coord, or
    	-- -   the modulus of the number pair formed from the new
    	--   X or Y coordinate and the other coordinate of this
    	--   vector that was not directly modified.

  SetXY (me: in out; Coord : XY)         raises ConstructionError  is static;
    	---C++:inline  
    	---Purpose:
    	-- Assigns:
    	-- -   the two coordinates of Coord to this unit vector,
	--   and then normalizes it.
    	-- Warning
    	-- Remember that all the coordinates of a unit vector are
    	-- implicitly modified when any single one is changed directly.
    	-- Exceptions
    	-- Standard_ConstructionError if either of the following
    	-- is less than or equal to gp::Resolution():
    	-- -   the modulus of Coord, or
    	-- -   the modulus of the number pair formed from the new
    	--   X or Y coordinate and the other coordinate of this
    	--   vector that was not directly modified.


  Coord (me; Index : Integer)   returns Real
    	---C++:inline  
        --- Purpose :
        --  For this unit vector returns the coordinate of range Index :
        --  Index = 1 => X is returned
        --  Index = 2 => Y is returned    
	-- Raises OutOfRange if Index != {1, 2}.
      raises OutOfRange
      is static;

  Coord (me; Xv, Yv : out Real) is static;
    	---C++:inline  
    	---Purpose: For this unit vector returns its two coordinates Xv and Yv.
	-- Raises OutOfRange if Index != {1, 2}.

  X (me)  returns Real          is static;
      	---C++:inline
    	--- Purpose: For this unit vector, returns its X coordinate.  
  Y (me)  returns Real          is static;
    	---C++:inline  
    	--- Purpose: For this unit vector, returns its Y coordinate.  

  XY (me)  returns XY           is static;
        ---C++: inline
        ---C++: return const& 
    	--- Purpose: For this unit vector, returns its two coordinates as a number pair.

        --- Purpose : Comparison between Directions
        --  The precision value is an input data.

  IsEqual (me; Other : Dir2d; AngularTolerance : Real)  returns Boolean
     is static;
       ---C++: inline     
       --- Purpose : 
       --  Returns True if the two vectors have the same direction 
       -- i.e. the angle between this unit vector and the
       -- unit vector Other is less than or equal to AngularTolerance.


  IsNormal (me; Other : Dir2d; AngularTolerance : Real)  returns Boolean
     is static;
        ---C++: inline     
        --- Purpose :
        --  Returns True if the angle between this unit vector and the
    	-- unit vector Other is equal to Pi/2 or -Pi/2 (normal)
    	-- i.e. Abs(Abs(<me>.Angle(Other)) - PI/2.) <= AngularTolerance


  IsOpposite (me; Other : Dir2d; AngularTolerance : Real)  returns Boolean
     is static;
        ---C++: inline     
        --- Purpose :
        --  Returns True if the angle between this unit vector and the
    	-- unit vector Other is equal to Pi or -Pi (opposite).
    	-- i.e.  PI - Abs(<me>.Angle(Other)) <= AngularTolerance


  IsParallel (me; Other : Dir2d; AngularTolerance : Real)  returns Boolean
     is static;
        ---C++: inline    
        --- Purpose :
        --  returns true if if the angle between this unit vector and unit
    	-- vector Other is equal to 0, Pi or -Pi.
    	-- i.e.  Abs(Angle(<me>, Other)) <= AngularTolerance or
    	--  PI - Abs(Angle(<me>, Other)) <= AngularTolerance

  Angle (me; Other : Dir2d)   returns Real   is static;
        --- Purpose :
        --  Computes the angular value in radians between <me> and 
        --  <Other>. Returns the angle in the range [-PI, PI].


  Crossed (me; Right : Dir2d)  returns Real  is static;
        ---C++: inline
        --- Purpose : 
        --  Computes the cross product between two directions.
        ---C++: alias operator ^


  Dot (me; Other : Dir2d)   returns Real   is static;
        ---C++: inline
        --- Purpose : Computes the scalar product
        ---C++: alias operator *




  Reverse (me : in out)         is static;
        ---C++: inline

  Reversed (me)  returns Dir2d  is static;
        ---C++: inline
    	---C++: alias operator -  
        --- Purpose : Reverses the orientation of a direction


  Mirror (me : in out; V : Dir2d)           is static;

  Mirrored (me; V : Dir2d)  returns Dir2d   is static;

        --- Purpose :
        --  Performs the symmetrical transformation of a direction
        --  with respect to the direction V which is the center of 
        --  the  symmetry.

  

  Mirror (me : in out; A : Ax2d)            is static;

  Mirrored (me; A : Ax2d)  returns Dir2d    is static;
      --- Purpose :
        --  Performs the symmetrical transformation of a direction
        --  with respect to an axis placement which is the axis
        --  of the symmetry.

  

  Rotate (me : in out; Ang : Real)          is static;
        ---C++: inline
	
  Rotated (me; Ang : Real)   returns Dir2d  is static;
	--- Purpose :
        --  Rotates a direction.  Ang is the angular value of 
        --  the rotation in radians.
        ---C++: inline

  Transform (me : in out; T : Trsf2d)          is static;

  Transformed (me; T : Trsf2d)  returns Dir2d  is static;
        ---C++: inline      

        --- Purpose :
        --  Transforms a direction with the "Trsf" T.
        --- Warnings :
        --  If the scale factor of the "Trsf" T is negative then the
        --  direction <me> is reversed.



fields

    coord : XY;

end;
