-- Created on: 2000-10-23
-- Created by: Pavel TELKOV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package XDEDRAW 

    ---Purpose: Provides DRAW commands for work with DECAF data structures

uses
    Draw

is

    class Shapes;
    	---Purpose: Provides functions for work with shapes and assemblies

    class Colors;
    	---Purpose: Provides functions for work with colors

    class Layers;
    	---Purpose: Provides functions for work with layers

    class Props;
    	---Purpose: Provides functions for work with geometric properties  
	
    class Common; 
    	---Purpose: Provides common commands for work XDE

    Init (di: in out Interpretor from Draw);
    	---Purpose: Initializes all the functions

    Factory (theDI : out Interpretor from Draw);
    ---Purpose: Loads all Draw commands of  TKXDEDRAW. Used for plugin.

end XDEDRAW;
