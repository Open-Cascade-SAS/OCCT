-- Created on: 1995-01-25
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class PresentationManager from PrsMgr
inherits TShared from MMgt

  ---Purpose: A framework to manage 3D displays, graphic entities and their updates.
  -- Used in the AIS package (Application Interactive Services), to enable the advanced user to define the
  -- default display mode of a new interactive object which extends the list of signatures and types.
  -- Definition of new display types is handled by calling the presentation algorithms provided by the StdPrs package.

uses 

  StructureManager    from Graphic3d,
  PresentableObject   from PrsMgr,
  ListOfPresentations from PrsMgr,
  Length,NameOfColor  from Quantity,
  Color               from Quantity,
  Transformation      from Geom,
  NameOfMaterial      from Graphic3d,
  Presentation        from PrsMgr,
  View                from V3d,
  ViewManager         from Visual3d,
  ShadingAspect       from Prs3d,
  Presentation        from Prs3d

raises

  NoSuchObject from Standard

is

  Create (theStructureManager : ViewManager from Visual3d)
  returns PresentationManager from PrsMgr;
  ---Purpose:
  -- Creates a framework to manage displays and graphic entities with the 3D view theStructureManager.

  Display (me           : mutable;
           thePrsObject : PresentableObject from PrsMgr;
           theMode      : Integer from Standard = 0)
  ---Purpose: Displays the presentation of the object in the given Presentation manager with the given mode.
  --          The mode should be enumerated by the object which inherits PresentableObject.
  is static;

  Erase (me           : mutable;
         thePrsObject : PresentableObject from PrsMgr;
         theMode      : Integer from Standard = 0)
  ---Level: public
  ---Purpose: erases the presentation of the object in the given
  --          Presentation manager with the given mode.
  is static;

  Clear (me           : mutable;
         thePrsObject : PresentableObject from PrsMgr;
         theMode      : Integer from Standard = 0)
  is virtual;
  ---Purpose:
  -- Clears the presentation of the presentable object thePrsObject in this framework with the display mode theMode.

  SetVisibility (me           : mutable;
                 thePrsObject : PresentableObject from PrsMgr;
                 theMode      : Integer from Standard;
                 theValue     : Boolean from Standard);
  ---Purpose: Sets the visibility of presentable object.

  Highlight (me           : mutable;
             thePrsObject : PresentableObject from PrsMgr;
             theMode      : Integer from Standard = 0)
  ---Purpose: Highlights the presentation of the presentable object
  -- thePrsObject in this framework with the display mode theMode.
  is static;

  Unhighlight (me           : mutable;
               thePrsObject : PresentableObject from PrsMgr;
               theMode      : Integer from Standard = 0)
  ---Purpose: Removes highlighting from the presentation of the
  -- presentable object thePrsObject in this framework with the display mode theMode.
  is static;

  SetDisplayPriority (me;
                      thePrsObject : PresentableObject from PrsMgr;
                      theMode      : Integer from Standard;
                      theNewPrior  : Integer from Standard);
  ---Purpose:
  -- Sets the display priority theNewPrior of the
  -- presentable object thePrsObject in this framework with the display mode theMode.

  DisplayPriority (me;
                   thePrsObject : PresentableObject from PrsMgr;
                   theMode      : Integer from Standard)
  returns Integer from Standard;
  ---Purpose:
  -- Returns the display priority of the presentable object
  -- thePrsObject in this framework with the display mode theMode.

  SetZLayer (me           : mutable;
             thePrsObject : PresentableObject from PrsMgr;
             theLayerId   : Integer from Standard)
  is static;
  ---Purpose: Set Z layer ID for all presentations of the object.

  GetZLayer (me;
             thePrsObject : PresentableObject from PrsMgr)
  returns Integer from Standard is static;
  ---Purpose: Get Z layer ID assigned to all presentations of the object.
  -- Method returns -1 value if object has no presentations and is
  -- impossible to get layer index.

  IsDisplayed (me;
               thePrsObject : PresentableObject from PrsMgr;
               theMode: Integer from Standard = 0)
  --Purpose: Returns true if the presentation of the presentable
  -- object thePrsObject in this framework with the display mode theMode is displayed.
  returns Boolean from Standard
  is static;

  IsHighlighted (me;
                 thePrsObject : PresentableObject from PrsMgr;
                 theMode: Integer from Standard = 0)
  ---Purpose: Returns true if the presentation of the presentable
  -- object thePrsObject in this framework with the display mode theMode is highlighted.
  returns Boolean from Standard
  is static;

  Update (me;
          thePrsObject : PresentableObject from PrsMgr;
          theMode      : Integer from Standard = 0)
  ---Purpose: Updates the presentation of the presentable object
  -- thePrsObject in this framework with the display mode theMode.
  is static;

---Category: Immediate display methods.

  BeginImmediateDraw (me : mutable);
  ---Purpose: Resets the transient list of presentations previously displayed in immediate mode
  -- and begins accumulation of new list by following AddToImmediateList()/Color()/Highlight() calls.

  ClearImmediateDraw (me : mutable);
  ---Purpose: Resets the transient list of presentations previously displayed in immediate mode.

  AddToImmediateList (me     : mutable;
                      thePrs : Presentation from Prs3d);
  ---Purpose: Stores thePrs in the transient list of presentations to be displayed in immediate mode.
  -- Will be taken in account in EndImmediateDraw method.

  EndImmediateDraw (me      : mutable;
                    theView : View from V3d);
  ---Purpose: Allows rapid drawing of the view theView by avoiding an update of the whole background.

  IsImmediateModeOn (me) returns Boolean from Standard;
  ---C++: inline
  ---Purpose: Returns true if Presentation Manager is accumulating transient list of presentations to be displayed in immediate mode.

---Category: Hilighting methods.

  Color (me           : mutable;
         thePrsObject : PresentableObject from PrsMgr;
         theColor     : NameOfColor from Quantity = Quantity_NOC_YELLOW;
         theMode      : Integer from Standard = 0;
         theSelObj    : PresentableObject from PrsMgr = NULL)
  ---Purpose: Highlights the graphic object thePrsObject in the color theColor.
  -- thePrsObject has the display mode theMode;
  -- this has the default value of 0, that is, the wireframe display mode.
  is static;

  BoundBox (me           : mutable;
            thePrsObject : PresentableObject from PrsMgr;
            theMode      : Integer from Standard = 0)
  ---Purpose: highlights the boundbox of the presentation
  is static;

---Category: references to other presentation.

  Connect (me             : mutable;
           thePrsObject   : PresentableObject from PrsMgr;
           theOtherObject : PresentableObject from PrsMgr;
           theMode        : Integer from Standard = 0;
           theOtherMode   : Integer from Standard = 0)
  is static;

---Category: Transformation methods.

  Transform (me                : mutable;
             thePrsObject      : PresentableObject from PrsMgr;
             theTransformation : Transformation from Geom;
             theMode           : Integer from Standard = 0)
  ---Purpose:
  -- Sets the transformation theTransformation for the presentable object thePrsObject.
  -- thePrsObject has the display mode theMode; this has the default value of 0, that is, the wireframe display mode.
  is static;

  StructureManager (me) returns StructureManager from Graphic3d
  is static;
  ---C++: inline
  ---C++: return const&
  ---Purpose: Returns the structure manager.

  SetShadingAspect (me           : mutable;
                    thePrsObject : PresentableObject from PrsMgr;
                    theColor     : NameOfColor from Quantity;
                    theMaterial  : NameOfMaterial from Graphic3d;
                    theMode      : Integer from Standard = 0)
  ---Purpose: this method will change the color and the aspect of the presentations containing shaded structures.
  is static;

  SetShadingAspect (me               : mutable;
                    thePrsObject     : PresentableObject from PrsMgr;
                    theShadingAspect : ShadingAspect from Prs3d;
                    theMode          : Integer from Standard = 0)
  ---Purpose: this method will change the color and the aspect of the presentations containing shaded structures.
  is static;

---Category: Private & deferred methods.

  HasPresentation (me;
                   thePrsObject : PresentableObject from PrsMgr;
                   theMode      : Integer from Standard = 0)
  returns Boolean from Standard
  is static;
  ---Purpose: Returns true if there is a presentation of the
  -- presentable object thePrsObject in this framework, thePrsObject having the display mode theMode.

  Presentation (me;
                thePrsObject : PresentableObject from PrsMgr;
                theMode      : Integer from Standard = 0;
                theToCreate  : Boolean from Standard = Standard_False;
                theSelObj    : PresentableObject from PrsMgr = NULL)
  returns Presentation from PrsMgr
  is static;
  ---Purpose: Returns the presentation Presentation of the presentable object thePrsObject in this framework.
  -- When theToCreate is true - automatically creates presentation for specified mode when not exist.
  -- Optional argument theSelObj specifies parent decomposed object to inherit its view affinity.

  RemovePresentation (me           : mutable;
                      thePrsObject : PresentableObject from PrsMgr;
                      theMode      : Integer from Standard = 0)
  returns Boolean from Standard
  ---Purpose: Removes a presentation of the presentable object thePrsObject to this framework. thePrsObject has the display mode theMode.
  is protected;

fields

  myStructureManager : ViewManager         from Visual3d  is protected;
  myImmediateModeOn  : Integer             from Standard  is protected;
  myImmediateList    : ListOfPresentations from PrsMgr    is protected;
  myImmediateView    : View                from V3d       is protected;
  mySelectionColor   : Color               from Quantity  is protected;

end PresentationManager from PrsMgr;
