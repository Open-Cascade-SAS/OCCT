-- Created on: 1997-09-11
-- Created by: Philippe MANGIN
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred class ElementaryCriterion from FEmTool inherits  TShared  from  MMgt

	---Purpose:  defined J Criteria to used in minimisation 

uses
   Vector  from  math, 
   Matrix  from  math,  
   HArray2OfReal  from  TColStd, 
   HArray2OfInteger  from TColStd 
    
raises 
  NotImplemented,   
  DomainError

is
    Set(me  :  mutable;   
        Coeff : HArray2OfReal) 
	 ---Purpose: Set the coefficient of the Element (the  Curve)
    is  static;
     
    Set(me : mutable; 
        FirstKnot  :  Real; 
        LastKnot   :  Real) 
	---Purpose: Set the definition interval of the Element         
    is virtual;  
     
    DependenceTable(me)  
    returns  HArray2OfInteger  from TColStd 
	---Purpose: To know if two dimension are independent.        
    is  deferred;  
    
    Value  (me  : mutable) 
    	---Purpose: To Compute J(E) where E  is the current Element        
    returns  Real  is  deferred;
     
    Hessian(me  :  mutable ;
	    Dim1  :  Integer; 
	    Dim2  :  Integer;
            H  :  out  Matrix  from  math) 
    ---Purpose: To Compute J(E)  the coefficients of Hessian matrix of
    --          J(E) wich are crossed derivatives in dimensions <Dim1>
    --          and  <Dim2>.          
     raises  DomainError -- If DependenceTable(Dimension1,Dimension2) is False 
     is  deferred;  
   
    Gradient(me   : mutable; 
	     Dim  :  Integer;
             G    :  out  Vector  from  math)     	 
    ---Purpose: To Compute the  coefficients in the dimension <dim> 
    --          of  the  J(E)'s  Gradient where E  is  the current  Element
    is  deferred;

fields 
  myCoeff           :  HArray2OfReal  is  protected; 
  myFirst,  myLast  :  Real is  protected;
end ElementaryCriterion;



