-- Created on: 2004-04-08
-- Created by: Sergey ZARITCHNY <szy@opencascade.com>
-- Copyright (c) 2004-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class NamedShapeDriver from BinMNaming inherits ADriver from BinMDF

	---Purpose: NamedShape  Attribute Driver.

uses
    SRelocationTable from BinObjMgt,
    RRelocationTable from BinObjMgt,
    Persistent       from BinObjMgt,
    MessageDriver    from CDM,
    Attribute        from TDF, 
    ShapeSet         from BinTools,
    LocationSet      from BinTools

is
    Create (theMessageDriver:MessageDriver from CDM)
        returns NamedShapeDriver from BinMNaming;

    NewEmpty (me)  returns Attribute from TDF;

    Paste(me; Source     : Persistent from BinObjMgt;
              Target     : Attribute from TDF;
              RelocTable : out RRelocationTable from BinObjMgt)
        returns Boolean from Standard;

    Paste(me; Source     : Attribute from TDF;
              Target     : in out Persistent from BinObjMgt;
              RelocTable : out SRelocationTable from BinObjMgt);
    
    ReadShapeSection (me: mutable; theIS: in out IStream from Standard);
      ---Purpose: Input the shapes from Bin Document file

    WriteShapeSection (me: mutable; theOS: in out OStream from Standard);
      ---Purpose: Output the shapes into Bin Document file

    Clear (me:mutable);
      ---Purpose: Clear myShapeSet 
       
    SetFormatNb(me: mutable; theFormat : Integer from Standard);  
    ---C++: inline 
    ---Purpose: set the format of topology  
    --          First : does not write CurveOnSurface UV Points into the file
    --                  on reading calls Check() method.
    --          Second: stores CurveOnSurface UV Points.

    GetFormatNb(me) returns Integer from Standard; 
    ---Purpose: get the format of topology  
    ---C++: inline 
    
    GetShapesLocations(me: mutable) returns LocationSet from BinTools; 
    ---Purpose: get the format of topology  
    ---C++: return &
    ---C++: inline 
    
fields
     
    myShapeSet          : ShapeSet from BinTools; 
    myFormatNb          : Integer  from Standard;
end NamedShapeDriver;
