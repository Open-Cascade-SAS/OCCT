-- Created on: 1996-10-11
-- Created by: Christian CAILLET
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SelectSubordinate  from IGESSelect  inherits SelectExtract

    ---Purpose : This selections uses Subordinate Status as sort criterium
    --           It is an integer number which can be :
    --           0 Independant
    --           1 Physically Dependant
    --           2 Logically Dependant
    --           3 Both (recorded)
    --           + to sort :
    --           4 : 1 or 3  ->  at least Physically
    --           5 : 2 or 3  ->  at least Logically
    --           6 : 1 or 2 or 3 -> any kind of dependance
    --             (corresponds to 0 reversed)

uses AsciiString from TCollection, Transient, InterfaceModel
 
is
 
    Create (status : Integer) returns mutable SelectSubordinate;
    ---Purpose : Creates a SelectSubordinate with a status to be sorted

    Status (me) returns Integer;
    ---Purpose : Returns the status used for sorting
 
    Sort (me; rank : Integer; ent : Transient; model : InterfaceModel)
        returns Boolean;
    ---Purpose : Returns True if <ent> is an IGES Entity with Subordinate
    --           Status matching the criterium

    ExtractLabel (me) returns AsciiString from TCollection;
    ---Purpose : Returns the Selection criterium : "IGES Entity, Independant"
    --           etc...

fields

    thestatus : Integer;

end SelectSubordinate;
