-- Created on: 2000-05-24
-- Created by: data exchange team
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Application from XCAFApp inherits Application from TDocStd

    ---Purpose: Implements an Application for the DECAF documents

uses
    SequenceOfExtendedString from TColStd,
    Document from TDocStd

is

    Create returns mutable Application from XCAFApp is protected;


    ---Purpose: methods from CDF_Application
    --          ============================


    Formats(me: mutable; Formats: out SequenceOfExtendedString from TColStd) 
    is redefined;    


    ResourcesName (me: mutable) returns CString from Standard is redefined;

    ---Purpose: methods from TDocStd_Application
    --          ================================

    InitDocument (me; aDoc : Document from TDocStd) is redefined;
    ---Purpose: Set XCAFDoc_DocumentTool attribute
    
    ---API: method for initialisation

    GetApplication (myclass) returns Application from XCAFApp;
    ---Purpose: Initializes (for the first time) and returns the 
    --          static object (XCAFApp_Application)
    --          This is the only valid method to get XCAFApp_Application
    --          object, and it should be called at least once before
    --          any actions with documents in order to init application

end Application;
