-- Created on: 1993-01-08
-- Created by: Philippe DAUTRY
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

deferred generic class Builder from Sweep(TheShape as any)
    

	---Purpose: This  is   a  signature class  describing services
	--          strictly required    by  the    Swept   Primitives
	--          algorithms, from the Topology Data Structure .
	--          


uses

    Orientation from TopAbs
is

    MakeCompound (me; aCompound : out TheShape)
    	---Purpose: Returns an empty Compound.
    is deferred;

    MakeCompSolid (me; aCompSolid : out TheShape)
    	---Purpose: Returns an empty CompSolid.
    is deferred;

    MakeSolid (me; aSolid : out TheShape)
    	---Purpose: Returns an empty Solid.
    is deferred;

    MakeShell (me; aShell : out TheShape)
    	---Purpose: Returns an empty Shell.
    is deferred;

    MakeWire (me; aWire : out TheShape)
    	---Purpose: Returns an empty Wire.
    is deferred;
    
    Add(me; aShape1 : in out TheShape; 
	    aShape2 : in     TheShape;
    	    Orient  : in     Orientation from TopAbs)
    	---Purpose: Adds the Shape 1 in the Shape 2, set to
    	--          <Orient> orientation.
    is deferred;
    
    Add(me; aShape1 : in out TheShape; 
	    aShape2 : in     TheShape)
    	---Purpose: Adds the Shape 1 in the Shape 2.
    is deferred;

end Builder from Sweep;


