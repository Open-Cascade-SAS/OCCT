-- Created on: 1994-11-30
-- Created by: Frederic MAUPAS
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Tool from TopoDSToStep

    ---Purpose: This Tool Class provides Information to build
    --          a ProSTEP Shape model from a Cas.Cad BRep.                 

uses

    Vertex from TopoDS,
    Edge   from TopoDS,
    Wire   from TopoDS,
    Face   from TopoDS,
    Shell  from TopoDS,
    Shape  from TopoDS,
    
    DataMapOfShapeTransient from MoniTool,
    
    TopologicalRepresentationItem from StepShape
    
is 

--  -----------------------------------------------------------
--  Constructor
--  -----------------------------------------------------------

    Create returns Tool from TopoDSToStep;
    
    Create(M : DataMapOfShapeTransient from MoniTool;
    	   FacetedContext : Boolean from Standard) 
    	returns Tool from TopoDSToStep;
    
    Init(me : in out;
    	 M : DataMapOfShapeTransient from MoniTool;
      	 FacetedContext : Boolean from Standard);

--  -----------------------------------------------------------
--  Fields update methods
--  -----------------------------------------------------------


    IsBound(me : in out;
    	    S  : Shape from TopoDS) 
    	returns Boolean from Standard;
	
    Bind(me : in out;
    	 S  : Shape from TopoDS;
	 T  : TopologicalRepresentationItem from StepShape);
	 
    Find(me : in out;
    	 S  : Shape from TopoDS)
    	returns TopologicalRepresentationItem from StepShape;

    Faceted(me) returns Boolean from Standard;

    SetCurrentShell(me : in out;
    	    	    S  : Shell from TopoDS);
		    
    CurrentShell(me) returns Shell from TopoDS;
    	---C++: return const &


    SetCurrentFace(me : in out;
    	    	   F  : Face from TopoDS);
		    
    CurrentFace(me) returns Face from TopoDS;
    	---C++: return const &


    SetCurrentWire(me : in out;
    	    	   W  : Wire from TopoDS);
		    
    CurrentWire(me) returns Wire from TopoDS;
    	---C++: return const &


    SetCurrentEdge(me : in out;
    	    	   E  : Edge from TopoDS);
		    
    CurrentEdge(me) returns Edge from TopoDS;
    	---C++: return const &


    SetCurrentVertex(me : in out;
    	    	     V  : Vertex from TopoDS);
		    
    CurrentVertex(me) returns Vertex from TopoDS;
    	---C++: return const &
    
    Lowest3DTolerance(me) returns Real from Standard;

    SetSurfaceReversed(me : in out;
    	    	       B  : Boolean from Standard);
		       
    SurfaceReversed(me) returns Boolean from Standard;

    Map (me) returns DataMapOfShapeTransient from MoniTool;
        ---C++: return const &

    PCurveMode (me) returns Integer;
    	---Purpose: Returns mode for writing pcurves
	--          (initialized by parameter write.surfacecurve.mode)
    
fields

    myDataMap         : DataMapOfShapeTransient from MoniTool;
    
    myFacetedContext  : Boolean from Standard;
    
    myLowestTol       : Real from Standard;
    
    myCurrentShell    : Shell from TopoDS;
    
    myCurrentFace     : Face from TopoDS;
    
    myCurrentWire     : Wire from TopoDS;
    
    myCurrentEdge     : Edge from TopoDS;
    
    myCurrentVertex   : Vertex from TopoDS;

    myReversedSurface : Boolean from Standard;
    
    myPCurveMode      : Integer from Standard;
    
end Tool;
