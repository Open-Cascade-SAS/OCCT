-- File:	StepShape_DimensionalLocation.cdl
-- Created:	Tue Apr 18 16:42:58 2000 
-- Author:	Andrey BETENEV
-- Generator:	ExpToCas (EXPRESS -> CASCADE/XSTEP Translator) V1.0
-- Copyright:	Matra Datavision 1999

class DimensionalLocation from StepShape
inherits ShapeAspectRelationship from StepRepr

    ---Purpose: Representation of STEP entity DimensionalLocation

uses
    HAsciiString from TCollection,
    ShapeAspect from StepRepr

is
    Create returns DimensionalLocation from StepShape;
	---Purpose: Empty constructor

end DimensionalLocation;
