-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.




class VectorOrDirection from StepGeom inherits SelectType from StepData

	-- <VectorOrDirection> is an EXPRESS Select Type construct translation.
	-- it gathers : Vector, Direction

uses

	Vector,
	Direction
is

	Create returns VectorOrDirection;
	---Purpose : Returns a VectorOrDirection SelectType

	CaseNum (me; ent : Transient) returns Integer;
	---Purpose: Recognizes a VectorOrDirection Kind Entity that is :
	--        1 -> Vector
	--        2 -> Direction
	--        0 else

	Vector (me) returns any Vector;
	---Purpose : returns Value as a Vector (Null if another type)

	Direction (me) returns any Direction;
	---Purpose : returns Value as a Direction (Null if another type)


end VectorOrDirection;

