-- Created on: 1995-12-01
-- Created by: EXPRESS->CDL V0.2 Translator
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class CompositeTextWithExtent from StepVisual 

inherits CompositeText from StepVisual 

uses

	PlanarExtent from StepVisual, 
	HAsciiString from TCollection, 
	HArray1OfTextOrCharacter from StepVisual
is

	Create returns mutable CompositeTextWithExtent;
	---Purpose: Returns a CompositeTextWithExtent


	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCollectedText : mutable HArray1OfTextOrCharacter from StepVisual) is redefined;

	Init (me : mutable;
	      aName : mutable HAsciiString from TCollection;
	      aCollectedText : mutable HArray1OfTextOrCharacter from StepVisual;
	      aExtent : mutable PlanarExtent from StepVisual) is virtual;

	-- Specific Methods for Field Data Access --

	SetExtent(me : mutable; aExtent : mutable PlanarExtent);
	Extent (me) returns mutable PlanarExtent;

fields

	extent : PlanarExtent from StepVisual;

end CompositeTextWithExtent;
