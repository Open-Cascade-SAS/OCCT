-- Created on: 1993-05-07
-- Created by: Jacques GOUSSARD
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class RstInt from IntPatch

    ---Purpose: trouver les points d intersection entre la ligne de
    --          cheminement et les arcs de restriction

uses Polygo     from IntPatch,
     Line       from IntPatch,
     HSurface   from Adaptor3d,
     TopolTool  from Adaptor3d

raises DomainError from Standard

is

    PutVertexOnLine(myclass;
                    L         : in out Line from IntPatch; 
                    Surf      : HSurface from Adaptor3d; 
                    Domain    : TopolTool from Adaptor3d; 
                    OtherSurf : HSurface from Adaptor3d; 
                    OnFirst   : Boolean from Standard ;
                    Tol       : Real from Standard;
                    hasBeenAdded: Boolean from Standard = Standard_False)

    	raises DomainError from Standard;
    	--- The exception is raised if the Line from is neither
    	--  a WLine nor a RLine.

end RstInt;
