-- Created on: 2002-10-31
-- Created by: Michael SAZONOV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class DocumentRetrievalDriver from BinLDrivers inherits RetrievalDriver from PCDM

uses
    HeaderData                  from Storage,
    Position                    from Storage,
    AsciiString                 from TCollection,
    ExtendedString              from TCollection,
    Document                    from PCDM,
    Document                    from CDM,
    Application                 from CDM,
    MessageDriver               from CDM,
    ADriverTable                from BinMDF,
    RRelocationTable            from BinObjMgt,
    Persistent                  from BinObjMgt,
    Label                       from TDF,
    IStream                     from Standard,
    MapOfInteger                from TColStd,
    DocumentSection             from BinLDrivers,
    VectorOfDocumentSection     from BinLDrivers

is
    -- ===== Public methods =====

    Create returns mutable DocumentRetrievalDriver from BinLDrivers;
        ---Purpose: Constructor

    SchemaName          (me)
        returns ExtendedString from TCollection is redefined virtual;
        ---Purpose: pure virtual method definition

    Make                (me : mutable; PD : Document from PCDM;
                                       TD : Document from CDM)
        is redefined virtual;
        ---Purpose: pure virtual method definition

    CreateDocument      (me : mutable)
        returns Document from CDM is redefined virtual;
        ---Purpose: pure virtual method definition

    Read(me:mutable; theFileName:    ExtendedString from TCollection;
                     theNewDocument: Document    from CDM;
                     theApplication: Application from CDM) is redefined virtual;
        ---Purpose: retrieves the content of the file into a new Document.

    AttributeDrivers  (me : mutable; theMsgDriver: MessageDriver from CDM)
        returns ADriverTable from BinMDF
        is virtual;

    -- ===== Protected methods =====

    ReadSubTree (me: mutable; theIS   : in out IStream from Standard;
                              theData : Label from TDF)
        returns Integer from Standard
        is virtual protected;
        ---Purpose: Read the tree from the stream <theIS> to <theLabel>

    ReadInfoSection(me: mutable; theFile : AsciiString from TCollection;
                                 theData : in out HeaderData from Storage)
        returns Position from Storage is protected;
        ---Purpose: Read the  info  section  of  theFile into theData,
        --          return a file  position  corresponding to the info
        --          section end
    
    ReadSection    (me: mutable;
                    theSection : in out DocumentSection from BinLDrivers;
                    theDoc     : Document    from CDM;
                    theIS      : in out IStream from Standard)
        is virtual protected; 
        ---Purpose: define the procedure of reading a section to file.

    ReadShapeSection (me: mutable;
                      theSection : in out DocumentSection from BinLDrivers;
                      theIS      : in out IStream from Standard; 
    	    	      isMess     : Boolean from Standard = Standard_False)
        is virtual protected; 
	
    CheckShapeSection (me: mutable;
                      thePos : Position from Storage;
                      theIS  : in out IStream from Standard)
        is virtual protected; 
	 
    PropagateDocumentVersion(me: mutable; theVersion : Integer from Standard) 
    	is virtual protected; 
	
    WriteMessage(me: mutable; theMessage : ExtendedString from TCollection)
        is protected;
        ---Purpose: write  theMessage  to  the  MessageDriver  of  the
        --          Application
    
fields
    -- use one self-increasing buffer for an attribute
    myPAtt      : Persistent            from BinObjMgt;
    myDrivers   : ADriverTable          from BinMDF    is protected;
    myRelocTable: RRelocationTable      from BinObjMgt is protected;
    myMsgDriver : MessageDriver         from CDM;
    -- map of type ID of attributes registered in file header but not having a driver
    myMapUnsupported :  MapOfInteger    from TColStd;

    mySections  : VectorOfDocumentSection from BinLDrivers;

end DocumentRetrievalDriver;
