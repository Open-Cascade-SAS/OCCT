-- Created on: 2000-10-31
-- Created by: Vladislav ROMASHKO
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class Common from QANewBRepNaming inherits BooleanOperationFeat from QANewBRepNaming

uses
 
    Label from TDF, 
    BooleanOperation from BRepAlgoAPI

is
 
    Create returns Common from QANewBRepNaming;

    Create(ResultLabel : Label from TDF) 
    returns Common from QANewBRepNaming;

    Load (me; MakeShape : in out BooleanOperation from BRepAlgoAPI);
  

end Cut;
