-- Created on: 1997-10-22
-- Created by: Jean-Louis Frenkel
-- Copyright (c) 1997-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

---Copy:	 Matra Datavision 1997

deferred class Application from CDM inherits Transient from Standard

uses Document           from CDM,
     MetaData           from CDM,
     Reference          from CDM,
     MessageDriver      from CDM,
     Manager            from Resource,
     ExtendedString     from TCollection
is

    Retrieve(me: mutable; aMetaData: MetaData from CDM; UseStorageConfiguration: Boolean from Standard)
    returns Document from CDM
    is deferred private;


    DocumentVersion(me: mutable; aMetaData: MetaData from CDM)
    returns Integer from Standard
    is deferred private;
    ---Purpose: returns -1 if the metadata has no modification counter.
    
    SetDocumentVersion(me; aDocument: Document from CDM; aMetaData: MetaData from CDM)
    is protected;

    SetReferenceCounter(me:mutable ; aDocument: Document from CDM; aReferenceCounter: Integer from Standard)
    is protected;
    
    Resources(me: mutable)
    returns Manager from Resource
    is deferred;
    ---Purpose: the manager returned by  this virtual  method will be
    --          used to search for Format`.Retrieval  resource items. 
    --          
    
    MessageDriver(me: mutable) returns MessageDriver from CDM
    is virtual;
    ---Purpose: By default returns a NullMessageDriver;

    BeginOfUpdate(me:mutable; aDocument: Document from CDM)
    is virtual;
    ---Purpose: this method is called before the update of a document.
    --         By default, writes in MessageDriver().

    EndOfUpdate(me:mutable; aDocument: Document from CDM; Status: Boolean from Standard; ErrorString: ExtendedString from TCollection)
    is virtual;
    ---Purpose: this method is called affter the update of a document.
    --         By default, writes in MessageDriver().

    Write(me: mutable; aString: ExtString from Standard);
    ---Purpose: writes the string in the application MessagerDriver.

friends     

    class Reference from CDM,
    class MetaData from CDM

end Application from CDM;
