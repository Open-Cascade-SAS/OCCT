-- File:        BrepWithVoids.cdl
-- Created:     Mon Dec  4 12:02:24 1995
-- Author:      EXPRESS->CDL V0.2 Translator
-- Copyright:   Matra-Datavision 1993




class RWBrepWithVoids from RWStepShape

	---Purpose : Read & Write Module for BrepWithVoids

uses Check from Interface,
     StepReaderData from StepData,
     StepWriter from StepData,
     BrepWithVoids from StepShape,
     EntityIterator from Interface,
     ShareTool from Interface

is

	Create returns RWBrepWithVoids;

	ReadStep (me; data : StepReaderData; num : Integer;
	              ach : in out Check; ent : mutable BrepWithVoids from StepShape);

	WriteStep (me; SW : in out StepWriter; ent : BrepWithVoids from StepShape);

	Share(me; ent : BrepWithVoids from StepShape; iter : in out EntityIterator);

    	Check(me; ent : BrepWithVoids from StepShape; shares : ShareTool; ach : in out Check);

end RWBrepWithVoids;
