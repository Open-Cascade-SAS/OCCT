-- Created on: 2000-10-20
-- Created by: Julia DOROVSKIKH
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class MidPointPresentation from DsgPrs

uses
    Presentation from Prs3d,
    Drawer       from Prs3d,
    Pnt   from gp,
    Lin   from gp,
    Circ  from gp,
    Elips from gp,
    Ax2   from gp

is
    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  theAxe       : Ax2 from gp;
		  MidPoint     : Pnt from gp;
	          Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
    	    	  first        : Boolean from Standard);
	           ---Purpose: draws the representation of a MidPoint between
	           --          two vertices.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  theAxe       : Ax2 from gp;
		  MidPoint     : Pnt from gp;
		  Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
	       	  Point1       : Pnt from gp;
		  Point2       : Pnt from gp;
    	    	  first        : Boolean from Standard);
		   ---Purpose: draws the representation of a MidPoint between
		   --          two lines or linear segments.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  aCircle      : Circ from gp;
		  MidPoint     : Pnt from gp;
		  Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
	       	  Point1       : Pnt from gp;
		  Point2       : Pnt from gp;
    	    	  first        : Boolean from Standard);
		   ---Purpose: draws the representation of a MidPoint between
		   --          two entire circles or two circular arcs.

    Add( myclass; aPresentation: Presentation from Prs3d;
    	    	  aDrawer      : Drawer from Prs3d;
		  anElips      : Elips from gp;
		  MidPoint     : Pnt from gp;
		  Position     : Pnt from gp;
	       	  AttachPoint  : Pnt from gp;
	       	  Point1       : Pnt from gp;
		  Point2       : Pnt from gp;
    	    	  first        : Boolean from Standard);
		   ---Purpose: draws the representation of a MidPoint between
		   --          two entire ellipses or two elliptic arcs.

end MidPointPresentation;
