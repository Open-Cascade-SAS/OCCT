-- Created on: 1999-05-13
-- Created by: data exchange team
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ConvertCurve3dToBezier from ShapeUpgrade inherits SplitCurve3d from ShapeUpgrade

    ---Purpose: converts/splits a 3d curve of any type to a list of beziers

uses

    HSequenceOfCurve from TColGeom,
    HSequenceOfReal from TColStd

is

    Create returns ConvertCurve3dToBezier from ShapeUpgrade;
    	---Purpose: Empty constructor
    
    SetLineMode(me:mutable; mode: Boolean);
    	---Purpose: Sets mode for conversion Geom_Line to bezier.
    	---C++: inline
    
    GetLineMode(me) returns Boolean;
    	---Purpose: Returns the Geom_Line conversion mode.
    	---C++: inline
    
    SetCircleMode(me:mutable; mode: Boolean);
    	---Purpose: Sets mode for conversion Geom_Circle to bezier.
    	---C++: inline
    
    GetCircleMode(me) returns Boolean;
    	---Purpose: Returns the Geom_Circle conversion mode.
    	---C++: inline
    
    SetConicMode(me:mutable; mode: Boolean);
    	---Purpose: Returns the Geom_Conic conversion mode.
    	---C++: inline
    
    GetConicMode(me) returns Boolean;
    	---Purpose: Performs converting and computes the resulting shape.
    	---C++: inline
    
    Compute(me: mutable) is redefined;
    	---Purpose: Converts curve into a list of beziers, and stores the 
    	--          splitting parameters on original curve.
    
    Build (me: mutable; Segment: Boolean) is redefined;
    	---Purpose: Splits a list of beziers computed by Compute method according
	--          the split values and splitting parameters.
    
    Segments(me) returns HSequenceOfCurve from TColGeom is private;
    	---Purpose: Returns the list of bezier curves correspondent to original
	--          curve.
    
    SplitParams(me) returns HSequenceOfReal from TColStd;
    	---Purpose: Returns the list of splitted parameters in original curve
	--          parametrisation.
    
fields

   mySegments   : HSequenceOfCurve from TColGeom;
   mySplitParams: HSequenceOfReal from TColStd;
   myLineMode   : Boolean;
   myCircleMode : Boolean;
   myConicMode  : Boolean;
    
end ConvertCurve2dToBezier;
 
