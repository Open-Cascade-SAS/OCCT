-- Created on: 2000-05-18
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package IntTools

 ---Purpose: Contains classes for intersection and classification
 ---         purposes and accompanying classes
uses
    
    TCollection, 
    TopoDS, 
    TopAbs, 
    TColStd, 
    BRepAdaptor, 
    BRepTopAdaptor,
    SortTools, 
    TopTools, 
    math,
    gp, 
    Bnd,
    Adaptor3d,
    GeomAdaptor,
    Geom,
    Geom2d,
    GeomInt,  
    GeomAbs,
    GeomAPI,
    Extrema,
    IntPatch, 
    IntSurf, 
    BRepClass3d, 
    TColgp, 
    MMgt, 
    Geom2dHatch, 
    
    BOPCol

is
    class Context; 
    class ShrunkRange; 
    --
    class Range;         
    class CommonPrt; 
    class Root; 
    class Compare; 
    class CompareRange;     

    class  EdgeEdge;

    class  EdgeFace;

    class  FClass2d;

    --class  LineConstructor;

    -----
    class MarkedRangeSet;

    class BaseRangeSample;

    class CurveRangeSample;

    class SurfaceRangeSample;

    class CurveRangeLocalizeData;

    class SurfaceRangeLocalizeData;

    class BeanFaceIntersector;


    class  Curve;

    class  PntOnFace;
    class  PntOn2Faces; 
      
    class  TopolTool;

    class  FaceFace;

    class  Tools; 

    generic class CArray1;   
    ---
    ---                 I  n  s  t  a  n  t  i  a  t  i  o  n  s  
    ---   
    imported SequenceOfPntOn2Faces; 
    --
    imported SequenceOfCurves; 
 
    
    imported SequenceOfRanges; 

    class  CArray1OfInteger  instantiates  
     CArray1(Integer from Standard); 
  
    class  CArray1OfReal  instantiates  
     CArray1(Real from Standard); 
  
    imported SequenceOfRoots; 
  
    imported Array1OfRoots;  
     
    imported Array1OfRange; 
  
    class  QuickSort         instantiates  
     QuickSort from SortTools   (Root from IntTools, 
                    Array1OfRoots from IntTools, 
                    Compare from IntTools); 
        
    class  QuickSortRange    instantiates  
     QuickSort from SortTools   (Range from IntTools, 
                    Array1OfRange from IntTools, 
                    CompareRange from IntTools); 
    imported SequenceOfCommonPrts;        
  
    imported IndexedDataMapOfTransientAddress; 
    

    imported ListOfCurveRangeSample;
    

    imported ListIteratorOfListOfCurveRangeSample;

    imported ListOfSurfaceRangeSample;

    imported ListIteratorOfListOfSurfaceRangeSample;

    imported ListOfBox;

    imported ListIteratorOfListOfBox;
 
    class CurveRangeSampleMapHasher;

    class SurfaceRangeSampleMapHasher;
    
    imported MapOfCurveSample;
    
    imported MapIteratorOfMapOfCurveSample;
        
    imported MapOfSurfaceSample;
        
    imported MapIteratorOfMapOfSurfaceSample;
    
    imported DataMapOfCurveSampleBox;
    
    imported DataMapIteratorOfDataMapOfCurveSampleBox;

    imported DataMapOfSurfaceSampleBox;

    imported DataMapIteratorOfDataMapOfSurfaceSampleBox;
    -----------------------------------------------------
    --  Block  of  static  functions  
    -----------------------------------------------------  
    Length  (E : Edge from TopoDS) 
     returns  Real  from  Standard; 
    ---Purpose:  returns the length of the edge;  

    RemoveIdenticalRoots  (aSeq  :out SequenceOfRoots from IntTools; 
                  anEpsT:    Real from Standard); 
    ---Purpose: Remove from  the  sequence aSeq the Roots  that  have  
    --          values ti and tj such as  |ti-tj]  <  anEpsT.     

    SortRoots (aSeq  :out SequenceOfRoots from IntTools; 
            anEpsT:    Real from Standard);  
    ---Purpose: Sort the sequence aSeq of the Roots to arrange the 
    --          Roons  in  increasing  order  
    
    FindRootStates  (aSeq  :out SequenceOfRoots from IntTools; 
                     anEpsNull:    Real from Standard);
    ---Purpose: Find the states (before  and  after) for  each  Root  
    --          from  the sequence aSeq 
     
    Parameter (P          : Pnt   from gp; 
                Curve      : Curve from Geom; 
                aParm      : out Real  from  Standard) 
        returns  Integer from Standard;          
 
    GetRadius(C:  Curve  from  BRepAdaptor; 
           t1,t3:Real  from  Standard; 
            R:out Real  from  Standard) 
        returns  Integer from Standard;    
  

    PrepareArgs(C:  in out Curve  from  BRepAdaptor;  
                tMax,tMin:  Real  from  Standard; 
                Discret  :  Integer from Standard;    
                Deflect  :  Real  from  Standard;  
                anArgs   :  out  CArray1OfReal  from IntTools) 
        returns  Integer from Standard; 

end IntTools; 



