-- Created on: 1995-03-28
-- Created by: Yves FRICAUD
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Substitution from BRepTools 

	---Purpose: A tool to substitute subshapes by other shapes.
	--          
    	--          
    	--          The user use the method Substitute to define the
    	--          modifications. 
    	--          A set of shapes is designated to replace a initial
    	--          shape. 
    	--
    	--          The method Build reconstructs a new Shape with the
    	--          modifications.The Shape and the new shape are 
    	--          registered.
    	--          

uses
    Shape                     from TopoDS,
    ListOfShape               from TopTools,	
    DataMapOfShapeListOfShape from TopTools
    
raises
    
    NoSuchObject from Standard
is
    
    Create returns Substitution from BRepTools;
    
    Clear ( me : in out)
    	---Purpose: Reset all the fields.
    is static;

    Substitute (me : in out; 
    	    	OldShape  : Shape from TopoDS;
    	    	NewShapes : ListOfShape from TopTools)
    	---Purpose: <Oldshape> will be replaced by <NewShapes>.
    	--          
    	--          <NewShapes> can be empty , in this case <OldShape>
    	--          will disparate from its ancestors.
    	--          
    	--          if an item of <NewShapes> is oriented FORWARD.
    	--          it will be oriented as <OldShape> in its ancestors.
    	--          else it will be reversed.
    is static;
    
    
    Build (me : in out; S : Shape from TopoDS)
	---Purpose: Build NewShape from <S> if its subshapes has modified.
	--          
	--          The methods <IsCopied> and <Copy> allows you to keep
	--          the resul of <Build>
    is static;	    
    
    IsCopied(me; S : Shape from TopoDS) returns Boolean
	---Purpose: Returns   True if <S> has   been  replaced .
    is static;
    
    Copy(me; S : Shape from TopoDS) returns ListOfShape from TopTools
	---Purpose: Returns the set of shapes  substitued to <S> .
	---C++: return const &
    raises
    	NoSuchObject from Standard -- if ! IsCopied(S)
    is static;
    
fields

    myMap    : DataMapOfShapeListOfShape from TopTools;
    
end Substitution;
