-- Created on: 1992-05-27
-- Created by: Remi LEQUETTE
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class TEdge from BRep inherits TEdge from TopoDS

	---Purpose: The TEdge from BRep is  inherited from  the  TEdge
	--          from TopoDS. It contains the geometric data.
	--          
	--          The TEdge contains :
	--           
	--           * A tolerance.
	--           
	--           * A same parameter flag.
	--           
	--           * A same range flag.
	--           
	--           * A Degenerated flag.
	--           
	--           *  A  list   of curve representation.

uses
    TShape                    from TopoDS,
    ListOfCurveRepresentation from BRep

is
    Create returns mutable TEdge from BRep;
	---Purpose: Creates an empty TEdge.
	
    Tolerance(me) returns Real
	---C++: inline
    is static;
    	
    Tolerance(me : mutable; T : Real)
	---C++: inline
    is static;
    
    UpdateTolerance(me : mutable; T : Real)
	---Purpose: Sets the tolerance  to the   max  of <T>  and  the
	--          current  tolerance.
	--          
	---C++: inline
    is static;
    
    SameParameter(me) returns Boolean
    is static;
    
    SameParameter(me : mutable; S : Boolean)
    is static;
    
    SameRange(me) returns Boolean
    is static;
    
    SameRange(me : mutable; S : Boolean)
    is static;
    
    Degenerated(me) returns Boolean
    is static;
    
    Degenerated(me : mutable; S : Boolean)
    is static;
    
    Curves(me) returns ListOfCurveRepresentation from BRep
	---C++: return const &
	---C++: inline
    is static;
    
    ChangeCurves(me : mutable) returns ListOfCurveRepresentation from BRep
	---C++: return &
	---C++: inline
    is static;
    
    EmptyCopy(me) returns mutable TShape from TopoDS;
	---Purpose: Returns a copy  of the  TShape  with no sub-shapes.
    
fields

    myTolerance     : Real;
    myFlags         : Integer;
    myCurves        : ListOfCurveRepresentation from BRep;

end TEdge;
