-- Created on: 1994-01-24
-- Created by: Gilles DEBARBOUILLE
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class BooleanParameter from Dynamic

inherits
    Parameter from Dynamic     
    
	---Purpose: This class describes a parameter with a boolean 
	--          as value.

uses

   CString from Standard,
   OStream from Standard

is

    Create(aparameter : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> as name.

    returns mutable BooleanParameter from Dynamic;
    
    Create(aparameter : CString from Standard; 
           avalue : Boolean from Standard) 

    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> and <avalue>
    --          respectively as name and value.

    returns mutable BooleanParameter from Dynamic;
    
    Create(aparameter , avalue : CString from Standard)
    
    ---Level: Advanced 
    
    ---Purpose: Creates a boolean parameter with <aparameter> as name 
    --          and <avalue> as value. <avalue> is a CString with two possible
    --          values which are : "Standard_True" and "Standard_False".

    returns mutable BooleanParameter from Dynamic;
    
    Value(me) returns Boolean from Standard
    
    ---Level: Public 
    
    ---Purpose: Returns the boolean value <thevalue>.
    
    is static;
    
    Value (me : mutable ; avalue : Boolean from Standard)
    
    ---Level: Advanced 
    
    --- Purpose: Sets the field <thevalue> with the boolean value <avalue>

    is static;
    
    Dump(me ; astream : in out OStream from Standard)
    
    ---Level: Internal 
    
    ---Purpose: Useful for debugging.
    
    is redefined;
    
fields

    thevalue : Boolean from Standard;

end BooleanParameter;
