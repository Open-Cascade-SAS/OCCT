-- Created on: 2006-08-07
-- Created by: Galina KULIKOVA
-- Copyright (c) 2006-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class SplitSurfaceArea from ShapeUpgrade inherits SplitSurface from ShapeUpgrade

	---Purpose:Split surface in the parametric space 
        -- in according specified number of splits on the 



is
    Create returns mutable SplitSurfaceArea from ShapeUpgrade; 
    	---Purpose: Empty constructor.
    
    NbParts(me: mutable) returns Integer;
    ---C++: inline
    ---C++: return &
    ---Purpose:Set number of split for surfaces
    
    Compute(me: mutable; Segment: Boolean = Standard_True) is redefined;
    
fields

myNbParts : Integer; -- number of splitting

end SplitSurfaceArea;
