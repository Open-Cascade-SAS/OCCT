-- Created on: 1994-11-16
-- Created by: Marie Jose MARTZ
-- Copyright (c) 1994-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

package GeomToIGES

--- Purpose: Creation des entites geometriques de IGES
--           a partir des entites de Geom .

uses Interface, IGESData, IGESBasic, IGESConvGeom, IGESGeom, IGESSolid, IGESToBRep,
     gp, Geom, Geom2d, GeomConvert, GeomLProp, TColStd, TopoDS, TopTools,
     Transfer, TransferBRep,  BRep, TCollection, ElCLib

is

-- classes du package

    class GeomCurve;
    class GeomEntity;
    class GeomPoint;
    class GeomSurface;
    class GeomVector;

end GeomToIGES;
