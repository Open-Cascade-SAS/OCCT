-- Created on: 1993-01-09
-- Created by: CKY / Contract Toubro-Larsen ( SIVA )
-- Copyright (c) 1993-1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and/or modify it under
-- the terms of the GNU Lesser General Public License version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class VertexList from IGESSolid  inherits IGESEntity

        ---Purpose: defines VertexList, Type <502> Form Number <1>
        --          in package IGESSolid
        --          A vertex is a point in R3. A vertex is the bound of an
        --          edge and can participate in the bounds of a face.
        --          It contains one or more vertices.

uses

        Pnt          from gp,
        XYZ          from gp,
        HArray1OfXYZ from TColgp

raises OutOfRange

is

        Create returns VertexList;

        -- Specific Methods pertaining to the class

        Init (me       : mutable; 
              vertices : HArray1OfXYZ);
        ---Purpose : This method is used to set the fields of the class
        --           VertexList
        --       - vertices : the vertices in the list

        NbVertices (me) returns Integer;
        ---Purpose : return the number of vertices in the list

        Vertex (me; num : Integer) returns Pnt
        raises OutOfRange;
        ---Purpose : returns the num'th vertex in the list
        -- raises exception if num  <= 0 or num > NbVertices()

fields

--
-- Class    : IGESSolid_VertexList
--
-- Purpose  : Declaration of variables specific to the definition
--            of the Class VertexList.
--
-- Reminder : A VertexList instance is defined by :
--            an array of vertex
--

        theVertices : HArray1OfXYZ;

end VertexList;
