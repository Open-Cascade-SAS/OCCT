-- Created on: 1992-12-15
-- Created by: Christian CAILLET
-- Copyright (c) 1992-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WorkSession  from IFSelect  inherits TShared

    ---Purpose : This class can be used to simply manage a process such as
    --           splitting a file, extracting a set of Entities ...           
    --           It allows to manage different types of Variables : Integer or
    --           Text Parameters, Selections, Dispatches, in addition to a
    --           ShareOut. To each of these variables, a unique Integer
    --           Identifier is attached. A Name can be attached too as desired.

uses CString, AsciiString from TCollection, HAsciiString from TCollection,
     Messenger from Message,
     SequenceOfHAsciiString from TColStd, HSequenceOfHAsciiString from TColStd,
     DictionaryOfInteger from Dico,
     Type, SequenceOfTransient  from TColStd, SequenceOfInteger  from TColStd,
     HSequenceOfInteger from TColStd,  HArray1OfInteger from TColStd,
     DictionaryOfTransient from Dico, IndexedDataMapOfTransientTransient,
     Transient,  HSequenceOfTransient from TColStd,
     InterfaceModel from Interface, EntityIterator from Interface,
     Protocol from Interface, HGraph from Interface, Graph from Interface,
     CheckIterator from Interface,  GTool from Interface,
     ShareOut, IntParam, Signature,  Selection,  Dispatch,   WorkLibrary,
     ModelCopier,  GeneralModifier,  Modifier,   Transformer,
     SelectionIterator,  PacketList, SignatureList,  SignCounter,
     ReturnStatus, RemainMode, PrintCount

raises DomainError

is

	-- --    General Management    -- --

    Create returns mutable WorkSession;
    ---Purpose : Creates a Work Session
    --           It provides default, empty ShareOut and ModelCopier, which can
    --           be replaced (if required, should be done just after creation).

    SetErrorHandle (me : mutable; hand : Boolean);
    ---Purpose : Changes the Error Handler status (by default, it is not set)

    ErrorHandle (me) returns Boolean;
    ---Purpose : Returns the Error Handler status

    ShareOut (me) returns mutable ShareOut;
    ---Purpose : Returns the ShareOut defined at creation time
    ---C++ : return const &

    SetShareOut (me : mutable; shareout : mutable ShareOut);
    ---Purpose : Sets a new ShareOut. Fills Items which its content
    --  Warning : data from the former ShareOut are lost
    
    SetModeStat(me : mutable; theMode : Boolean);
    ---Purpose : Set value of mode responsible for precence of selections after loading
    -- If mode set to true that different selections will be accessible after loading
    -- else selections will be not accessible after loading( for economy memory in applicatios) 
    
    GetModeStat(me)  returns Boolean from Standard;
    ---Purpose : Return value of mode defining of filling selection during loading


    SetLibrary (me : mutable; lib : WorkLibrary);
    ---Purpose : Sets a WorkLibrary, which will be used to Read and Write Files

    WorkLibrary (me) returns WorkLibrary;
    ---Purpose : Returns the WorkLibrary. Null Handle if not yet set
    -- should be C++ : return const &

    SetProtocol (me : mutable; protocol : Protocol from Interface);
    ---Purpose : Sets a Protocol, which will be used to determine Graphs, to
    --           Read and to Write Files

    Protocol (me) returns Protocol;
    ---Purpose : Returns the Protocol. Null Handle if not yet set
    -- should be C++ : return const &

    SetSignType (me : mutable; signtype : Signature);
    ---Purpose : Sets a specific Signature to be the SignType, i.e. the
    --           Signature which will determine TypeName from the Model
    --           (basic function). It is recorded in the GTool
    --           This Signature is also set as "xst-sign-type" (reserved name)
    --           

    SignType    (me) returns Signature;
    ---Purpose : Returns the current SignType


    HasModel (me) returns Boolean;
    ---Purpose : Returns True is a Model has been set

    SetModel (me : mutable; model : InterfaceModel;
    	      clearpointed : Boolean = Standard_True);
    ---Purpose : Sets a Model as input : this will be the Model from which the
    --           ShareOut will work
    --           if <clearpointed> is True (default) all SelectPointed items
    --              are cleared, else they must be managed by the caller
    --           Remark : SetModel clears the Graph, recomputes it if a
    --           Protocol is set and if the Model is not empty, of course

    Model (me) returns InterfaceModel;
    ---Purpose : Returns the Model of the Work Session (Null Handle if none)
    -- should be C++ : return const &

    SetLoadedFile (me : mutable; filename : CString);
    ---Purpose : Stores the filename used for read for setting the model
    --           It is cleared by SetModel and ClearData(1)

    LoadedFile (me) returns CString;
    ---Purpose : Returns the filename used to load current model
    --           empty if unknown

    ReadFile (me : mutable; filename : CString) returns ReturnStatus;
    ---Purpose : Reads a file with the WorkLibrary (sets Model and LoadedFile)
    --           Returns a integer status which can be :
    --           RetDone if OK,  RetVoid if no Protocol not defined,
    --           RetError for file not found, RetFail if fail during read

    NbStartingEntities (me) returns Integer;
    ---Purpose : Returns the count of Entities stored in the Model, or 0

    StartingEntity (me; num : Integer) returns Transient;
    ---Purpose : Returns an  Entity stored in the Model of the WorkSession
    --           (Null Handle is no Model or num out of range)

    StartingNumber (me; ent : Transient) returns Integer;
    ---Purpose : Returns the Number of an Entity in the Model
    --           (0 if no Model set or <ent> not in the Model)

    NumberFromLabel (me; val : CString; afternum : Integer= 0) returns Integer;
    ---Purpose : From a given label in Model, returns the corresponding number
    --           Starts from first entity by Default, may start after a given
    --           number : this number may be given negative, its absolute value
    --           is then considered. Hence a loop on NumberFromLabel may be
    --           programmed (stop test is : returned value positive or null)
    --           
    --           Returns 0 if not found, < 0 if more than one found (first
    --           found in negative).
    --           If <val> just gives an integer value, returns it

    EntityLabel (me; ent : Transient) returns HAsciiString from TCollection;
    ---Purpose : Returns the label for <ent>, as the Model does
    --           If <ent> is not in the Model or if no Model is loaded, a Null
    --           Handle is returned

    EntityName     (me; ent : Transient) returns HAsciiString from TCollection;
    ---Purpose : Returns the Name of an Entity
    --           This Name is computed by the general service Name
    --           Returns a Null Handle if fails

    CategoryNumber (me; ent : Transient) returns Integer;
    ---Purpose : Returns the Category Number determined for an entity
    --           it is computed by the class Category
    --           An unknown entity (number 0) gives a value -1

    CategoryName   (me; ent : Transient) returns CString;
    ---Purpose : Returns the Category Name determined for an entity
    --           it is computed by the class Category
    --           Remark : an unknown entity gives an empty string

    ValidityName   (me; ent : Transient) returns CString;
    ---Purpose : Returns the Validity Name determined for an entity
    --           it is computed by the class SignValidity
    --           Remark : an unknown entity gives an empty string

    ClearData (me : mutable; mode : Integer)  is virtual;
    ---Purpose : Clears recorded data (not the items) according mode :
    --           1 : all Data : Model, Graph, CheckList, + ClearData 4
    --           2 : Graph and CheckList (they will then be recomputed later)
    --           3 : CheckList (it will be recomputed by ComputeCheck)
    --           4 : just content of SelectPointed and Counters
    --           Plus 0 : does nothing but called by SetModel
    --           ClearData is virtual, hence it can be redefined to clear
    --             other data of a specialised Work Session

    ComputeGraph (me : mutable; enforce : Boolean = Standard_False) returns Boolean;
    ---Purpose : Computes the Graph used for Selections, Displays ...
    --           If a HGraph is already set, with same model as given by method
    --           Model, does nothing. Else, computes a new Graph.
    --           If <enforce> is given True, computes a new Graph anyway.
    --           Remark that a call to ClearGraph will cause ComputeGraph to
    --           really compute a new Graph
    --           Returns True if Graph is OK, False else (i.e. if no Protocol
    --           is set, or if Model is absent or empty).

    HGraph (me : mutable) returns HGraph;
    ---Purpose : Returns the Computed Graph as HGraph (Null Handle if not set)

    Graph (me : mutable) returns Graph
    ---Purpose : Returns the Computed Graph, for Read only
        raises DomainError;
    --           Error if the Graph is not available
    ---C++ : return const &

    Shareds  (me : mutable; ent : Transient) returns HSequenceOfTransient;
    ---Purpose : Returns the list of entities shared by <ent> (can be empty)
    --           Returns a null Handle if <ent> is unknown

    Sharings (me : mutable; ent : Transient) returns HSequenceOfTransient;
    ---Purpose : Returns the list of entities sharing <ent> (can be empty)
    --           Returns a null Handle if <ent> is unknown

    IsLoaded (me) returns Boolean;
    ---Purpose : Returns True if a Model is defined and really loaded (not
    --           empty), a Protocol is set and a Graph has been computed.
    --           In this case, the WorkSession can start to work

    ComputeCheck (me : mutable; enforce : Boolean = Standard_False)
    	returns Boolean;
    ---Purpose : Computes the CheckList for the Model currently loaded
    --           It can then be used for displays, querries ...
    --           Returns True if OK, False else (i.e. no Protocol set, or Model
    --           absent). If <enforce> is False, works only if not already done
    --           or if a new Model has been loaded from last call.
    -- Remark : computation is enforced by every call to
    --          SetModel or RunTransformer

    ModelCheckList (me : mutable; complete : Boolean = Standard_True)
    	returns CheckIterator;
    ---Purpose : Returns the Check List for the Model currently loaded :
    --           <complete> = True  : complete (syntactic & semantic messages),
    --               computed if not yet done
    --           <complete> = False : only syntactic (check file form)

    CheckOne (me : mutable; ent : Transient; complete : Boolean = Standard_True)
    	returns CheckIterator;
    ---Purpose : Returns a Check for a single entity, under the form of a
    --           CheckIterator (this gives only one form for the user)
    --           if <ent> is Null or equates the current Model, it gives the
    --           Global Check, else the Check for the given entity
    --           <complete> as for ModelCheckList

    LastRunCheckList (me) returns CheckIterator;
    ---Purpose : Returns the Check List produced by the last execution of
    --           either : EvaluateFile(for Split), SendSplit, SendAll,
    --           SendSelected, RunTransformer-RunModifier
    --           Cleared by SetModel or ClearData(1)
    --           The field is protected, hence a specialized WorkSession may
    --           fill it

    	-- --    General Management on  Items (and Names)    -- --

    MaxIdent (me) returns Integer;
    ---Purpose : Returns the Maximum Value for an Item Identifier. It can be
    --           greater to the count of known Items, because some can have
    --           been removed

    Item (me; id : Integer) returns mutable Transient;
    ---Purpose : Returns an Item, given its Ident. Returns a Null Handle if
    --           no Item corresponds to this Ident.

    ItemIdent (me; item : Transient) returns Integer;
    ---Purpose : Returns the Ident attached to an Item in the WorkSession, or
    --           Zero if it is unknown

    NamedItem (me; name : CString) returns mutable Transient;
    ---Purpose : Returns the Item which corresponds to a Variable, given its
    --           Name (whatever the type of this Item).
    --           Returns a Null Handle if this Name is not recorded

    NamedItem (me; name : HAsciiString from TCollection) returns mutable Transient;
    ---Purpose : Same as above, but <name> is given through a Handle
    --           Especially Usefull with methods SelectionNames, etc...

    NameIdent (me; name : CString) returns Integer;
    ---Purpose : Returns the Ident attached to a Name, 0 if name not recorded

    HasName (me; item : Transient) returns Boolean;
    ---Purpose : Returns True if an Item of the WorkSession has an attached Name

    Name (me; item : Transient) returns HAsciiString from TCollection;
    ---Purpose : Returns the Name attached to an Item as a Variable of this
    --           WorkSession. If <item> is Null or not recorded, returns an
    --           empty string.

    AddItem (me : mutable; item : mutable Transient;
    	 active : Boolean = Standard_True)  returns Integer;
    ---Purpose : Adds an Item and returns its attached Ident. Does nothing
    --           if <item> is already recorded (and returns its attached Ident)
    --           <active> if True commands call to SetActive (see below)
    --           Remark : the determined Ident is used if <item> is a Dispatch,
    --           to fill the ShareOut

    AddNamedItem (me : mutable; name : CString; item : mutable Transient;
    	active : Boolean = Standard_True)  returns Integer;
    ---Purpose : Adds an Item with an attached Name. If the Name is already
    --           known in the WorkSession, the older item losts it
    --           Returns Ident if Done, 0 else, i.e. if <item> is null
    --           If <name> is empty, works as AddItem (i.e. with no name)
    --           If <item> is already known but with no attached Name, this
    --           method tries to attached a Name to it
    --           <active> if True commands call to SetActive (see below)

    SetActive (me : mutable; item : mutable Transient; mode : Boolean)
    	returns Boolean;
    ---Purpose : Following the type of <item> :
    --           - Dispatch : Adds or Removes it in the ShareOut & FileNaming
    --           - GeneralModifier : Adds or Removes it for final sending
    --             (i.e. in the ModelCopier)
    --           Returns True if it did something, False else (state unchanged)

    RemoveNamedItem (me : mutable; name : CString) returns Boolean;
    ---Purpose : Removes an Item from the Session, given its Name
    --           Returns True if Done, False else (Name not recorded)
    --           (Applies only on Item which are Named)

    RemoveName (me : mutable; name : CString) returns Boolean;
    ---Purpose : Removes a Name without removing the Item
    --           Returns True if Done, False else (Name not recorded)

    RemoveItem (me : mutable; item : Transient) returns Boolean;
    ---Purpose : Removes an Item given its Ident. Returns False if <id> is
    --           attached to no Item in the WorkSession. For a Named Item,
    --           also removes its Name.

    ClearItems (me : mutable);
    ---Purpose : Clears all the recorded Items : Selections, Dispatches,
    --           Modifiers, and Strings & IntParams, with their Idents & Names.
    --           Remark that if a Model has been loaded, it is not cleared.

    ItemLabel (me; id : Integer) returns HAsciiString from TCollection;
    ---Purpose : Returns a Label which illustrates the content of an Item,
    --           given its Ident. This Label is :
    --           - for a Text Parameter, "Text:<text value>"
    --           - for an Integer Parameter, "Integer:<integer value>"
    --           - for a Selection, a Dispatch or a Modifier, its Label
    --             (see these classes)
    --           - for any other kind of Variable, its cdl type

    ItemIdents (me; type : Type) returns HSequenceOfInteger from TColStd;
    ---Purpose : Fills a Sequence with the List of Idents attached to the Items
    --           of which Type complies with (IsKind) <type> (alphabetic order)
    --           Remark : <type> = TYPE(Standard_Transient) gives all the
    --           Idents which are suitable in the WorkSession

    ItemNames (me; type : Type) returns HSequenceOfHAsciiString from TColStd;
    ---Purpose : Fills a Sequence with the list of the Names attached to Items
    --           of which Type complies with (IsKind) <type> (alphabetic order)
    --           Remark : <type> = TYPE(Standard_Transient) gives all the Names

    ItemNamesForLabel (me; label : CString) returns HSequenceOfHAsciiString;
    ---Purpose : Fills a Sequence with the NAMES of the control items, of which
    --           the label matches <label> (contain it) : see NextIdentForLabel
    --           Search mode is fixed to "contained"
    --           If <label> is empty, returns all Names

    NextIdentForLabel (me; label : CString; id : Integer; mode : Integer = 0)
    	returns Integer;
    ---Purpose : For query by Label with possible iterations
    --           Searches the Ident of which Item has a Label which matches a
    --           given one, the search starts from an initial Ident.
    --           Returns the first found Ident which follows <id>, or ZERO
    --           
    --           The search must start with <id> = 0, it returns the next Ident
    --           which matches. To iterate, call again this method which this
    --           returned value as <id>. Once an Ident has been returned, the
    --           Item can be obtained by the method Item
    --           
    --           <mode> precises the required matching mode :
    --           - 0 (Default) : <label> must match exactly with the Item Label
    --           - 1 : <label> must match the exact beginning (the end is free)
    --           - 2 : <label> must be at least once wherever in the Item Label
    --           - other values are ignored

	-- --    List of Parameters    -- --
	-- They are Integer (IntParam) and Text (HAsciiString from TCollection)

    NewParamFromStatic (me : mutable; statname : CString; name : CString = "")
    	returns mutable Transient;
    ---Purpose : Creates a parameter as being bound to a Static
    --           If the Static is Integer, this creates an IntParam bound to
    --           it by its name. Else this creates a String which is the value
    --           of the Static.
    --           Returns a null handle if <statname> is unknown as a Static

    IntParam (me; id : Integer) returns mutable IntParam;
    ---Purpose : Returns an IntParam, given its Ident in the Session
    --           Null result if <id> is not suitable for an IntParam
    --           (undefined, or defined for another kind of variable)

    IntValue (me; it : IntParam) returns Integer;
    ---Purpose : Returns Integer Value of an IntParam

    NewIntParam (me : mutable; name : CString = "") returns mutable IntParam;
    ---Purpose : Creates a new IntParam. A Name can be set (Optional)
    --           Returns the created IntParam, or a Null Handle in case of
    --           Failure (see AddItem/AddNamedItem)

    SetIntValue (me : mutable; it : mutable IntParam; val : Integer)
    	returns Boolean;
    ---Purpose : Changes the Integer Value of an IntParam
    --           Returns True if Done, False if <it> is not in the WorkSession


    TextParam (me; id : Integer) returns mutable HAsciiString from TCollection;
    ---Purpose : Returns a TextParam, given its Ident in the Session
    --           Null result if <id> is not suitable for a TextParam
    --           (undefined, or defined for another kind of variable)

    TextValue (me; par : HAsciiString from TCollection)
    	 returns AsciiString from TCollection;
    ---Purpose : Returns Text Value of a TextParam (a String)
    --           or an empty string if <it> is not in the WorkSession

    NewTextParam (me : mutable; name : CString = "")
    	 returns mutable HAsciiString from TCollection;
    ---Purpose : Creates a new (empty) TextParam. A Name can be set (Optional)
    --           Returns the created TextParam (as an HAsciiString), or a Null
    --           Handle in case of Failure (see AddItem/AddNamedItem)

    SetTextValue (me : mutable; par : mutable HAsciiString from TCollection;
    	    	  val : CString)  returns Boolean;
    ---Purpose : Changes the Text Value of a TextParam (an HAsciiString)
    --           Returns True if Done, False if <it> is not in the WorkSession

	-- --    List of Signatures    -- --

    Signature (me; id : Integer) returns mutable Signature;
    ---Purpose : Returns a Signature, given its Ident in the Session
    --           Null result if <id> is not suitable for a Signature
    --           (undefined, or defined for another kind of variable)

    SignValue (me; sign : Signature; ent : Transient) returns CString;
    ---Purpose : Returns the Value computed by a Signature for an Entity
    --           Returns an empty string if the entity does not belong to the
    --           loaded model

	-- --    List of Selections    -- --

    Selection (me; id : Integer) returns mutable Selection;
    ---Purpose : Returns a Selection, given its Ident in the Session
    --           Null result if <id> is not suitable for a Selection
    --           (undefined, or defined for another kind of variable)

    EvalSelection (me; sel : Selection) returns EntityIterator
    ---Purpose : Evaluates the effect of a Selection applied on the input Model
    --           Returned Result remains empty if no input Model has been set
    	raises DomainError;
    --           If ErrorHandle has been set and if an Error occurs, the
    --           exception is caught and the result is returned empty
    --           Else, the exception remains raised

    Sources (me; sel : Selection) returns SelectionIterator;
    ---Purpose : Returns the Selections which are source of Selection, given
    --           its rank in the List of Selections (see SelectionIterator)
    --           Returned value is empty if <num> is out of range or if
    --           <sel> is not in the WorkSession

    SelectionResult (me; sel : Selection) returns
    	HSequenceOfTransient from TColStd  raises DomainError;
    ---Purpose : Returns the result of a Selection, computed by EvalSelection
    --           (see above) under the form of a HSequence (hence, it can be
    --           used by a frontal-engine logic). It can be empty
    --           Returns a Null Handle if <sel> is not in the WorkSession

    SelectionResultFromList (me; sel : Selection; list : HSequenceOfTransient)
    	returns  HSequenceOfTransient from TColStd  raises DomainError;
    ---Purpose : Returns the result of a Selection, by forcing its input with
    --           a given list <list> (unless <list> is Null).
    --               RULES :
    --           <list> applies only for a SelectDeduct kind Selection :
    --           its Input is considered : if it is a SelectDeduct kind
    --            Selection, its Input is considered, etc... until an Input
    --           is not a Deduct/Extract : its result is replaced by <list>
    --           and all the chain of deductions is applied


    SetItemSelection (me : mutable; item : mutable Transient;
    	    	    	   sel : mutable Selection)  returns Boolean;
    ---Purpose : Sets a Selection as input for an item, according its type :
    --           if <item> is a Dispatch : as Final Selection
    --           if <item> is a GeneralModifier (i.e. any kind of Modifier) :
    --             as Selection used to filter entities to modify
    --           <sel>  Null  causes this Selection to be nullified
    --           Returns False if <item> is not of a suitable type, or
    --             <item> or <sel> is not in the WorkSession

    ResetItemSelection (me : mutable; item : mutable Transient) returns Boolean;
    ---Purpose : Resets input Selection which was set by SetItemSelection
    --           Same conditions as for SetItemSelection
    --           Returns True if done, False if <item> is not in the WorkSession

    ItemSelection (me; item : Transient) returns mutable Selection;
    ---Purpose : Returns the Selection of a Dispatch or a GeneralModifier.
    --           Returns a Null Handle if none is defined or <item> not good type

	-- --    Counters    -- --
	-- a Counter can be used directly
	-- it can also be recorded as control item of the WorkSession, then :
	-- - it is cleared by ClearData (1 or 4)
	-- - when it is defined by a Selection, it can be recomputed

    SignCounter (me; id : Integer) returns mutable SignCounter;
    ---Purpose : Returns a SignCounter from its ident in the Session
    --           Null result if <id> is not suitable for a SignCounter
    --           (undefined, or defined for another kind of variable)

    ComputeCounter (me : mutable; counter : SignCounter;
    	    	    forced : Boolean=Standard_False)  returns Boolean;
    ---Purpose : Computes the content of a SignCounter when it is defined with
    --           a Selection, then returns True
    --           Returns False if the SignCounter is not defined with a
    --           Selection, or if its Selection Mode is inhibited
    --           <forced> to work around optimisations

    ComputeCounterFromList (me : mutable; counter : SignCounter;
    	    	list : HSequenceOfTransient; clear : Boolean = Standard_True)
    	    	    returns Boolean;
    ---Purpose : Computes the content of a SignCounter from an input list
    --           If <list> is Null, uses internal definition of the Counter :
    --             a Selection, else the whole Model (recomputation forced)
    --           If <clear> is True (D), starts from scratch
    --           Else, cumulates computations

	-- --    Dispatches (stored by ShareOut)    -- --

    AppliedDispatches (me) returns HSequenceOfInteger from TColStd;
    ---Purpose : Returns the ordered list of dispatches stored by the ShareOut

    ClearShareOut (me : mutable; onlydisp : Boolean);
    ---Purpose : Clears the list of Dispatches recorded by the ShareOut
    --           if <only> disp is True, tha's all. Else, clears also the lists
    --           of Modifiers recorded by the ShareOut

    Dispatch (me; id : Integer) returns mutable Dispatch;
    ---Purpose : Returns a Dispatch, given its Ident in the Session
    --           Null result if <id> is not suitable for a Dispatch
    --           (undefined, or defined for another kind of variable)


    DispatchRank (me; disp : Dispatch) returns Integer;
    ---Purpose : Returns the rank of a Dispatch in the ShareOut, or 0 if <disp>
    --           is not in the ShareOut or not in the WorkSession

    	-- --    Modifiers (cf also ModelCopier)    -- --
    	--   A Modifier can be applied to : final sending (all dispatches),
    	--   final sending but for one specific Dispatch, or another action
    	--   
    	--   Modifiers can be, either active for final sending to file (managed
    	--   by the ModelCopier), or not.
    	--   Here, Management of Modifiers (except the global list) concerns
    	--   only active Modifiers for the final sending.
    	--   But Criteria (Selection,Dispatch) are suitable for every kind of
    	--   Modifier, i.e. for GeneralModifier (also applies to IFAdapt kinds
    	--   of Modifiers, which apply during the Copy operation itself)

    ModelCopier (me) returns mutable ModelCopier;
    ---Purpose : Gives access to the complete ModelCopier

    SetModelCopier (me : mutable; copier : mutable ModelCopier);
    ---Purpose : Sets a new ModelCopier. Fills Items which its content
    ---Warning : all data recorded in the former ModelCopier are lost
    --           (thus, Final Modifiers become inactive)

    NbFinalModifiers (me; formodel : Boolean) returns Integer;
    ---Purpose : Returns the count of Modifiers applied to final sending
    --           Model Modifiers if <formodel> is True, File Modifiers else
    --           (i.e. Modifiers which apply once the Models have been filled)

    FinalModifierIdents (me; formodel : Boolean)
    	 returns HSequenceOfInteger from TColStd;
    ---Purpose : Fills a Sequence with a list of Idents, those attached to
    --           the Modifiers applied to final sending.
    --           Model Modifiers if <formodel> is True, File Modifiers else
    --           This list is given in the order in which they will be applied
    --           (which takes into account the Changes to Modifier Ranks)

    GeneralModifier (me; id : Integer)
    	returns mutable GeneralModifier;
    ---Purpose : Returns a Modifier, given its Ident in the Session
    --           Null result if <id> is not suitable for a Modifier
    --           (undefined, or defined for another kind of variable)

    ModelModifier (me; id : Integer) returns mutable Modifier;
    ---Purpose : Returns a Model Modifier, given its Ident in the Session,
    --           i.e. typed as a Modifier (not simply a GeneralModifier)
    --           Null result if <id> is not suitable for a Modifier
    --           (undefined, or defined for another kind of variable)

    ModifierRank (me; item : GeneralModifier) returns Integer;
    ---Purpose : Returns the Rank of a Modifier given its Ident. Model or File
    --           Modifier according its type (ModelModifier or not)
    --           Remember that Modifiers are applied sequencially following
    --           their Rank : first Model Modifiers then File Modifiers
    --           Rank is given by rank of call to AddItem and can be
    --           changed by ChangeModifierRank

    ChangeModifierRank (me : mutable;
    	formodel : Boolean; before, after : Integer) returns Boolean;
    ---Purpose : Changes the Rank of a Modifier in the Session :
    --           Model Modifiers if <formodel> is True, File Modifiers else
    --           the Modifier n0 <before> is put to n0 <after>
    --           Return True if Done, False if <before> or <after> out of range

    ClearFinalModifiers (me : mutable);
    ---Purpose : Removes all the Modifiers active in the ModelCopier : they
    --           become inactive and they are removed from the Session

    SetAppliedModifier (me : mutable; modif : mutable GeneralModifier;
    	    	        item : mutable Transient) returns Boolean;
    ---Purpose : Sets a GeneralModifier to be applied to an item :
    --           - item = ShareOut : applies for final sending (all dispatches)
    --           - item is a Dispatch : applies for this dispatch only
    --           Returns True if done, False if <modif> or <item> not in <me>

    ResetAppliedModifier (me : mutable; modif : mutable GeneralModifier)
    	returns Boolean;
    ---Purpose : Resets a GeneralModifier to be applied
    --           Returns True if done, False if <modif> was not applied

    UsesAppliedModifier (me; modif : GeneralModifier) returns mutable Transient;
    ---Purpose : Returns the item on which a GeneralModifier is applied :
    --           the ShareOut, or a given Dispatch
    --           Returns a Null Handle if <modif> is not applied

    	-- --    Transformation (without sending)    -- --

    Transformer (me; id : Integer) returns mutable Transformer;
    ---Purpose : Returns a Transformer, given its Ident in the Session
    --           Null result if <id> is not suitable for a Transformer
    --           (undefined, or defined for another kind of variable)

    RunTransformer (me : mutable; transf : Transformer)  returns Integer;
    ---Purpose : Runs a Transformer on starting Model, which can then be edited
    --           or replaced by a new one. The Protocol can also be changed.
    --           Fills LastRunCheckList
    --           
    --           Returned status is 0 if nothing done (<transf> or model
    --             undefined), positive if OK, negative else :
    --           0  : Nothing done
    --           1  : OK, edition on the spot with no change to the graph
    --                of dependances (purely local)
    --           2  : OK, model edited on the spot (graph recomputed, may
    --               have changed), protocol unchanged
    --           3  : OK, new model produced, same protocol
    --           4  : OK, model edited on the spot (graph recomputed),
    --                but protocol has changed
    --           5  : OK, new model produced, protocol has changed
    --           -1 : Error on the spot (slight changes), data may be corrupted
    --                (remark : corruption should not be profound)
    --           -2 : Error on edition the spot, data may be corrupted
    --                (checking them is recommanded)
    --           -3 : Error with a new data set, transformation ignored
    --           -4 : OK as 4, but graph of dependances count not be recomputed
    --                (the former one is kept) : check the protocol

    RunModifier (me : mutable; modif : Modifier; copy : Boolean) 
    	returns Integer;
    ---Purpose : Runs a Modifier on Starting Model. It can modify entities, or
    --           add new ones. But the Model or the Protocol is unchanged.
    --           The Modifier is applied on each entity of the Model. See also
    --             RunModifierSelected
    --           Fills LastRunCheckList
    --           
    --           <copy> : if True, a new data set is produced which brings
    --             the modifications (Model + its Entities)
    --           if False, data are modified on the spot
    --           
    --           It works through a TransformStandard defined with <modif>
    --           Returned status as RunTransformer : 0 nothing done, >0 OK,
    --           <0 problem, but only between -3 and 3 (protocol unchanged)
    --           Remark : <copy> True will give <effect> = 3 or -3

    RunModifierSelected  (me : mutable; modif : Modifier;
    	sel : Selection;  copy : Boolean) 
    	returns Integer;
    ---Purpose : Acts as RunModifier, but the Modifier is applied on the list
    --           determined by a Selection, rather than on the whole Model
    --           If the selection is a null handle, the whole model is taken

    NewTransformStandard (me : mutable; copy : Boolean; name : CString = "")
    	 returns mutable Transformer;
    ---Purpose : Creates and returns a TransformStandard, empty, with its
    --           Copy Option (True = Copy, False = On the Spot) and an
    --           optional name.
    --           To a TransformStandard, the method SetAppliedModifier applies

    SetModelContent (me : mutable; sel : Selection; keep : Boolean)
    	returns Boolean;
    ---Purpose : Defines a new content from the former one
    --           If <keep> is True, it is given by entities selected by
    --              Selection <sel>  (and all shared entities)
    --           Else, it is given by all the former content but entities
    --              selected by the Selection <sel> (and properly shared ones)
    --           Returns True if done. Returns False if the selected list
    --           (from <sel>) is empty, hence nothing is done

	-- --    File and Transfer Management    -- --

    FilePrefix (me) returns HAsciiString from TCollection;
    ---Purpose : Returns the defined File Prefix. Null Handle if not defined

    DefaultFileRoot (me) returns HAsciiString from TCollection;
    ---Purpose : Returns the defined Default File Root. It is used for
    --           Dispatches which have no specific root attached.
    --           Null Handle if not defined

    FileExtension (me) returns HAsciiString from TCollection;
    ---Purpose : Returns the defined File Extension. Null Handle if not defined

    FileRoot (me; disp : Dispatch) returns HAsciiString from TCollection;
    ---Purpose : Returns the File Root defined for a Dispatch. Null if no
    --           Root Name is defined for it (hence, no File will be produced)

    SetFilePrefix (me : mutable; name : CString);
    ---Purpose : Defines a File Prefix

    SetDefaultFileRoot (me : mutable; name : CString) returns Boolean;
    ---Purpose : Defines a Default File Root Name. Clears it is <name> = ""
    --           Returns True if OK, False if <name> already set for a Dispatch

    SetFileExtension (me : mutable; name : CString);
    ---Purpose : Defines a File Extension

    SetFileRoot (me : mutable; disp : Dispatch; name : CString) returns Boolean;
    ---Purpose : Defines a Root for a Dispatch
    --           If <name> is empty, clears Root Name
    --           This has as effect to inhibit the production of File by <disp>
    --           Returns False if <disp> is not in the WorkSession or if a
    --           root name is already defined for it

    GiveFileRoot (me; file : CString) returns CString;
    ---Purpose : Extracts File Root Name from a given complete file name
    --           (uses OSD_Path)

    GiveFileComplete (me; file : CString) returns CString;
    ---Purpose : Completes a file name as required, with Prefix and Extension
    --           (if defined; for a non-defined item, completes nothing)

    ClearFile (me : mutable);
    ---Purpose : Erases all stored data from the File Evaluation
    --           (i.e. ALL former naming informations are lost)

    EvaluateFile (me : mutable);
    ---Purpose : Performs and stores a File Evaluation. The Results are a List
    --           of produced Models and a List of names (Strings), in parallel
    --           Fills LastRunCheckList

    NbFiles   (me) returns Integer;
    ---Purpose : Returns the count of produced Models

    FileModel (me; num : Integer) returns mutable InterfaceModel;
    ---Purpose : Returns a Model, given its rank in the Evaluation List

    FileName  (me; num : Integer) returns AsciiString from TCollection;
    ---Purpose : Returns the name of a file corresponding to a produced Model,
    --           given its rank in the Evaluation List

    BeginSentFiles (me : mutable; record : Boolean);
    ---Purpose : Commands file sending to clear the list of already sent files,
    --           commands to record a new one if <record> is True
    --           This list is managed by the ModelCopier when SendSplit is called
    --           It allows a global exploitation of the set of sent files

    SentFiles (me) returns HSequenceOfHAsciiString;
    ---Purpose : Returns the list of recorded sent files, or a Null Handle is
    --           recording has not been enabled


    SendSplit (me : mutable) returns Boolean;
    ---Purpose : Performs creation of derived files from the input Model
    --           Takes its data (sub-models and names), from result EvaluateFile
    --           if active, else by dynamic Evaluation (not stored)
    --           After SendSplit, result of EvaluateFile is Cleared
    --           Fills LastRunCheckList
    --           
    --           Works with the WorkLibrary which acts on specific type of Model
    --           and can work with File Modifiers (managed by the Model Copier)
    --           and a ModelCopier, which can work with Model Modifiers
    --           Returns False if, either WorkLibrary has failed on at least
    --           one sub-file, or the Work Session is badly conditionned
    --           (no Model defined, or FileNaming not in phase with ShareOut)

    EvalSplit (me) returns PacketList;
    ---Purpose : Returns an Evaluation of the whole ShareOut definition : i.e.
    --           how the entities of the starting model are forecast to be sent
    --           to various files :  list of packets according the dispatches,
    --           effective lists of roots for each packet (which determine the
    --           content of the corresponding file); plus evaluation of which
    --           entities are : forgotten (sent into no file), duplicated (sent
    --           into more than one file), sent into a given file.
    --           See the class PacketList for more details.

    SentList (me; count : Integer = -1)  returns EntityIterator;
    ---Purpose : Returns the list of Entities sent in files, accourding the
    --           count of files each one has been sent (these counts are reset
    --           by SetModel or SetRemaining(Forget) ) stored in Graph Status
    --           <count> = -1 (default) is for ENtities sent at least once
    --           <count> = 0 is for the Remaining List (entities not yet sent)
    --           <count> = 1 is for entities sent in one and only one file
    --             (the ideal case)
    --           Remaining Data are computed on each Sending/Copying output
    --           files (see methods EvaluateFile and SendSplit)
    --           Graph Status is 0 for Remaining Entity, <count> for Sent into
    --           <count> files
    --           This status is set to 0 (not yet sent) for all by SetModel
    --           and by SetRemaining(mode=Forget,Display)

    MaxSendingCount (me) returns Integer;
    ---Purpose : Returns the greater count of different files in which any of
    --           the starting entities could be sent.
    --           Before any file output, this count is 0.
    --           Ideal count is 1. More than 1 means that duplications occur.

    SetRemaining (me : mutable; mode : RemainMode) returns Boolean;
    ---Purpose : Processes Remaining data (after having sent files), mode :
    --           Forget  : forget remaining info (i.e. clear all "Sent" status)
    --           Compute : compute and keep remaining (does nothing if :
    --                 remaining is empty or if no files has been sent)
    --           Display : display entities recorded as remaining
    --           Undo    : restore former state of data (after Remaining(1) )
    --           Returns True if OK, False else (i.e. mode = 2 and Remaining
    --           List is either empty or takes all the entities, or mode = 3
    --           and no former computation of remaining data was done)


    SendAll (me : mutable; filename : CString;
    	     computegraph : Boolean = Standard_False) returns ReturnStatus;
    ---Purpose : Sends the starting Model into one file, without splitting,
    --           managing remaining data or anything else.
    --           <computegraph> true commands the Graph to be recomputed before
    --           sending : required when a Model is filled in several steps
    --           
    --           The Model and File Modifiers recorded to be applied on sending
    --           files are.
    --           Returns a status of execution : 
    --             Done if OK, 
    --             Void if no data available,
    --             Error if errors occured (work library is not defined), errors 
    --             during translation
    --             Fail if exception during translation is raised
    --             Stop if no disk space or disk, file is write protected
    --           Fills LastRunCheckList

    SendSelected (me : mutable; filename : CString; sel : Selection;
    	     computegraph : Boolean = Standard_False) returns ReturnStatus;
    ---Purpose : Sends a part of the starting Model into one file, without
    --           splitting. But remaining data are managed.
    --           <computegraph> true commands the Graph to be recomputed before
    --           sending : required when a Model is filled in several steps
    --           
    --           The Model and File Modifiers recorded to be applied on sending
    --           files are.
    --           Returns a status : Done if OK,  Fail if error during send,
    --            Error : WorkLibrary not defined, Void : selection list empty
    --           Fills LastRunCheckList

    WriteFile    (me : mutable; filename : CString) returns ReturnStatus;
    ---Purpose : Writes the current Interface Model globally to a File, and
    --           returns a write status which can be :
    --             Done OK, Fail file could not be written, Error no norm is selected
    -- Remark  : It is a simple, one-file writing, other operations are
    --           available (such as splitting ...) which calls SendAll

    WriteFile    (me : mutable; filename : CString; sel : Selection from IFSelect)
    	 returns ReturnStatus;
    ---Purpose : Writes a sub-part of the current Interface Model to a File,
    --           as defined by a Selection <sel>, recomputes the Graph, and
    --           returns a write status which can be :
    --             Done OK, Fail file could not be written, Error no norm is selected
    -- Remark  : It is a simple, one-file writing, other operations are
    --           available (such as splitting ...) which calls SendSelected

	-- --    Some General Purpose Selections    -- --

    NbSources (me; sel : Selection) returns Integer;
    ---Purpose : Returns the count of Input Selections known for a Selection,
    --           or 0 if <sel> not in the WorkSession. This count is one for a
    --           SelectDeduct / SelectExtract kind, two for SelectControl kind,
    --           variable for a SelectCombine (Union/Intersection), zero else

    Source (me; sel : Selection; num : Integer = 1) returns mutable Selection;
    ---Purpose : Returns the <num>th Input Selection of a Selection
    --           (see NbSources).
    --           Returns a Null Handle if <sel> is not in the WorkSession or if
    --           <num> is out of the range <1-NbSources>
    --           To obtain more details, see the method Sources

    IsReversedSelectExtract (me; sel : Selection) returns Boolean;
    ---Purpose : Returns True if <sel> a Reversed SelectExtract, False else

    ToggleSelectExtract (me : mutable; sel : mutable Selection) returns Boolean;
    ---Purpose : Toggles the Sense (Direct <-> Reversed) of a SelectExtract
    --           Returns True if Done, False if <sel> is not a SelectExtract or
    --           is not in the WorkSession

    SetInputSelection (me : mutable; sel, input : mutable Selection)
    	returns Boolean;
    ---Purpose : Sets an Input Selection (as <input>) to a SelectExtract or
    --           a SelectDeduct (as <sel>).
    --           Returns True if Done, False if <sel> is neither a
    --           SelectExtract nor a SelectDeduct, or not in the WorkSession


    SetControl (me : mutable; sel, sc : mutable Selection;
       	        formain : Boolean = Standard_True) returns Boolean;
    ---Purpose : Sets an Input Selection, Main if <formain> is True, Second else
    --           (as <sc>) to a SelectControl (as <sel>). Returns True if Done,
    --           False if <sel> is not a SelectControl, or <sc> or <sel> is not
    --           in the WorkSession

    CombineAdd  (me : mutable; selcomb, seladd : mutable Selection;
    	    	 atnum : Integer = 0)  returns Integer;
    ---Purpose : Adds an input selection to a SelectCombine (Union or Inters.).
    --           Returns new count of inputs for this SelectCombine if Done or
    --           0 if <sel> is not kind of SelectCombine, or if <seladd> or
    --           <sel> is not in the WorkSession
    --           By default, adding is done at the end of the list
    --           Else, it is an insertion to rank <atnum> (usefull for Un-ReDo)

    CombineRemove (me : mutable; selcomb, selrem : mutable Selection)
    	returns Boolean;
    ---Purpose : Removes an input selection from a SelectCombine (Union or
    --           Intersection). Returns True if done, False if <selcomb> is not
    --           kind of SelectCombine or <selrem> is not source of <selcomb>

    NewSelectPointed (me : mutable; list : HSequenceOfTransient; name : CString)
    	returns mutable Selection;
    ---Purpose : Creates a new Selection, of type SelectPointed, its content
    --           starts with <list>. A name must be given (can be empty)

    SetSelectPointed (me; sel : mutable Selection; list : HSequenceOfTransient;
    	    	      mode : Integer) returns Boolean;
    ---Purpose : Changes the content of a Selection of type SelectPointed
    --           According <mode> : 0  set <list> as new content (clear former)
    --             1  : adds <list> to actual content
    --            -1  : removes <list> from actual content
    --           Returns True if done, False if <sel> is not a SelectPointed

	-- --    Various Evaluations   -- --

    GiveSelection (me; selname : CString) returns Selection;
    ---Purpose : Returns a Selection from a Name :
    --           - the name of a Selection : this Selection
    --           - the name of a Signature + criteria between (..) : a new
    --             Selection from this Signature
    --           - an entity or a list of entities : a new SelectPointed
    --           Else, returns a Null Handle

    GiveList (me; obj : Transient) returns HSequenceOfTransient;
    ---Purpose : Determines a list of entities from an object :
    --           <obj> already HSequenceOfTransient : returned itself
    --           <obj> Selection : its Result of Evaluation is returned
    --           <obj> an entity of the Model : a HSequence which contains it
    --           else, an empty HSequence
    --           <obj> the Model it self : ALL its content (not only the roots)

    GiveList (me; first : CString; second : CString = "")
    	returns HSequenceOfTransient;
    ---Purpose : Computes a List of entities from two alphanums,
    --           first and second, as follows :
    --           if <first> is a Number or Label of an entity : this entity
    --           if <first> is a list of Numbers/Labels : the list of entities
    --           if <first> is the name of a Selection in <WS>, and <second>
    --             not defined, the standard result of this Selection
    --           else, let's consider "first second" : this whole phrase is
    --           splitted by blanks, as follows (RECURSIVE CALL) :
    --           - the leftest term is the final selection
    --           - the other terms define the result of the selection
    --           - and so on (the "leftest minus one" is a selection, of which
    --             the input is given by the remaining ...)

    GiveListFromList (me; selname : CString; ent : Transient)
    	returns HSequenceOfTransient;
    ---Purpose : Computes a List of entities from the model as follows
    --           <first> beeing a Selection or a combination of Selections,
    --             <ent> beeing an entity or a list
    --           of entities (as a HSequenceOfTransient) :
    --             the standard result of this selection applied to this list
    --           if <ent> is Null, the standard definition of the selection is
    --             used (which contains a default input selection)
    --           if <selname> is erroneous, a null handle is returned
    --           
    --           REMARK : selname is processed as <first second> of preceeding
    --             GiveList

    GiveListCombined (me; l1, l2 : HSequenceOfTransient; mode : Integer)
    	returns HSequenceOfTransient;
    ---Purpose : Combines two lists and returns the result, according to mode :
    --           <mode> < 0 : entities in <l1> AND NOT in <l2>
    --           <mode> = 0 : entities in <l1> AND in <l2>
    --           <mode> > 0 : entities in <l1> OR  in <l2>

    QueryCheckList (me : mutable; chl : CheckIterator);
    ---Purpose : Loads data from a check iterator to query status on it

    QueryCheckStatus (me; ent : Transient) returns Integer;
    ---Purpose : Determines check status for an entity regarding last call to
    --           QueryCheckList :
    --           -1 : <ent> unknown in the model, ignored
    --            0 : no check at all, immediate or inherited thru Graph
    --            1 : immediate warning (no fail), no inherited check
    --            2 : immediate fail, no inherited check
    --           +10 : idem but some inherited warning (no fail)
    --           +20 : idem but some inherited fail

    QueryParent (me; entdad, entson : Transient) returns Integer;
    ---Purpose : Determines if <entdad> is parent of <entson> (in the graph),
    --           returns : -1 if no; 0 if <entdad> = <entson>
    --           1 if immediate parent, > 1 if parent, gives count of steps

	-- --    Dumps, Evaluations (displayed on standard output)   -- --

    SetParams (me : mutable;
    	       params  : SequenceOfTransient;
    	       uselist : SequenceOfInteger);
    ---Purpose : Sets a list of Parameters, i.e. TypedValue, to be handled
    --           through an Editor
    --           The two lists are parallel, if <params> is longer than <uses>,
    --           surnumeral parameters are for general use
    --           
    --           EditForms are created to handle these parameters (list, edit)
    --           on the basis of a ParamEditor  xst-params-edit
    --           
    --           A use number dispatches the parameter to a given EditForm
    --           EditForms are defined as follows
    --           Name                Use   Means
    --           xst-params          all   All Parameters (complete list)
    --           xst-params-general  1     Generals
    --           xst-params-load     2     LoadFile (no Transfer)
    --           xst-params-send     3     SendFile (Write, no Transfer)
    --           xst-params-split    4     Split
    --           xst-param-read      5     Transfer on Reading
    --           xst-param-write     6     Transfer on Writing

    TraceStatics    (me; use : Integer; mode : Integer = 0);
    ---Purpose : Traces the Statics attached to a given use number
    --           If <use> is given positive (normal), the trace is embedded
    --           with a header and a trailer
    --           If <use> is negative, just values are printed
    --             (this allows to make compositions)
    --           Remark : use number  5 commands use -2 to be traced
    --           Remark : use numbers 4 and 6 command use -3 to be traced

    DumpShare (me);
    ---Purpose : Dumps contents of the ShareOut (on "cout")

    ListItems (me; label : CString = "");
    ---Purpose : Lists the Labels of all Items of the WorkSession
    --           If <label> is defined, lists labels which contain it

    ListFinalModifiers (me; formodel : Boolean);
    ---Purpose : Lists the Modifiers of the session (for each one, displays
    --           its Label). Listing is done following Ranks (Modifiers are
    --           invoked following their ranks)
    --           Model Modifiers if <formodel> is True, File Modifiers else

    DumpSelection (me; sel : Selection);
    ---Purpose : Lists a Selection and its Sources (see SelectionIterator),
    --           given its rank in the list

    DumpModel (me : mutable; level : Integer; S : Messenger from Message);
    ---Purpose : Lists the content of the Input Model (if there is one)
    --           According level : 0 -> gives only count of Entities and Roots
    --           1 -> Lists also Roots;  2 -> Lists all Entities (by TraceType)
    --           3 -> Performs a call to CheckList (Fails) and lists the result
    --           4 -> as 3 but all CheckList (Fails + Warnings)
    --           5,6,7  : as 3 but resp. Count,List,Labels by Fail
    --           8,9,10 : as 4 but resp. Count,List,Labels by message

    TraceDumpModel (me : mutable; mode : Integer);
    ---Purpose : Dumps the current Model (as inherited DumpModel), on currently
    --           defined Default Trace File (default is standard output)

    DumpEntity (me; ent : Transient; level : Integer; S : Messenger from Message);
    ---Purpose : Dumps a starting entity according to the current norm.
    --           To do this, it calls DumpEntity from WorkLibrary.
    --           <level> is to be interpreted for each norm : see specific
    --           classes of WorkLibrary for it. Generally, 0 if for very basic
    --           (only type ...), greater values give more and more details.

    PrintEntityStatus (me : mutable; ent : Transient; S : Messenger from Message);
    ---Purpose : Prints main informations about an entity : its number, type,
    --           validity (and checks if any), category, shareds and sharings..
    --           mutable because it can recompute checks as necessary

    TraceDumpEntity (me; ent : Transient; level : Integer);
    ---Purpose : Dumps an entity from the current Model as inherited DumpEntity
    --           on currently defined Default Trace File
    --           (<level> interpreted according to the Norm, see WorkLibrary)

    PrintCheckList (me; checklist : CheckIterator;
                    failsonly : Boolean; mode : PrintCount);
    ---Purpose : Prints a CheckIterator to the current Trace File, controlled
    --           with the current Model
    --           complete or fails only, according to <failsonly>
    --           <mode> defines the mode of printing
    --           0 : sequential, according entities; else with a CheckCounter
    --           1 : according messages, count of entities
    --           2 : id but with list of entities, designated by their numbers
    --           3 : as 2 but with labels of entities

    PrintSignatureList (me; signlist : SignatureList; mode : PrintCount);
    ---Purpose : Prints a SignatureList to the current Trace File, controlled
    --           with the current Model
    --           <mode> defines the mode of printing (see SignatureList)


    EvaluateSelection (me; sel : Selection);
    ---Purpose : Displays the list of Entities selected by a Selection (i.e.
    --           the result of EvalSelection).

    EvaluateDispatch (me; disp : Dispatch; mode : Integer = 0);
    ---Purpose : Displays the result of applying a Dispatch on the input Model
    --           (also shows Remainder if there is)
    --           <mode> = 0 (default), displays nothing else
    --           <mode> = 1 : displays also duplicated entities (because of
    --              this dispatch)
    --           <mode> = 2 : displays the entities of the starting Model
    --              which are not taken by this dispatch (forgotten entities)
    --           <mode> = 3 : displays both duplicated and forgotten entities
    --           Remark : EvaluateComplete displays these data evaluated for
    --           for all the dispatches, if there are several

    EvaluateComplete (me; mode : Integer = 0);
    ---Purpose : Displays the effect of applying the ShareOut on the input
    --           Model.
    --           <mode> = 0 (default) : displays only roots for each packet,
    --           <mode> = 1 : displays all entities for each packet, plus
    --             duplicated entities
    --           <mode> = 2 : same as <mode> = 1, plus displays forgotten
    --             entities (which are in no packet at all)

    ListEntities (me; iter : EntityIterator; mode : Integer);
    ---Purpose : Internal method which displays an EntityIterator
    --           <mode> 0 gives short display (only entity numbers)
    --           1 gives a more complete trace (1 line per Entity)
    --           (can be used each time a trace has to be output from a list)
    --           2 gives a form suitable for givelist : (n1,n2,n3...)

fields

    theerrhand   : Boolean;
    theshareout  : ShareOut;

    thelibrary   : WorkLibrary;
    theprotocol  : Protocol from Interface;
    themodel     : InterfaceModel;
    thegraph     : HGraph     is protected;
    theloaded    : AsciiString;
    thegtool     : GTool from Interface;

    thecheckdone : Boolean;
    thechecklist : CheckIterator;
    thecheckrun  : CheckIterator  is protected;  -- (LastRunCheckList)
    thecheckana  : AsciiString;

    theitems     : IndexedDataMapOfTransientTransient  is protected;
    thenames     : DictionaryOfTransient    is protected;

    thecopier    : ModelCopier;    -- produces + memorizes transferred data
    theoldel     : InterfaceModel;
	themodelstat : Boolean;
end WorkSession;
