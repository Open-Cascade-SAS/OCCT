-- Created on: 1999-05-11
-- Created by: Sergei ZERTCHANINOV
-- Copyright (c) 1999 Matra Datavision
-- Copyright (c) 1999-2014 OPEN CASCADE SAS
--
-- This file is part of Open CASCADE Technology software library.
--
-- This library is free software; you can redistribute it and / or modify it
-- under the terms of the GNU Lesser General Public version 2.1 as published
-- by the Free Software Foundation, with special exception defined in the file
-- OCCT_LGPL_EXCEPTION.txt. Consult the file LICENSE_LGPL_21.txt included in OCCT
-- distribution for complete text of the license and disclaimer of any warranty.
--
-- Alternatively, this file may be used under the terms of Open CASCADE
-- commercial license or contractual agreement.

class EdgeConnect  from ShapeFix

    ---Purpose : Makes vertices to be shared to connect edges,
    --           updates positions and tolerances for shared vertices.
    --           Accepts edges bounded by two vertices each.

uses 
    DataMapOfShapeShape from TopTools,
    DataMapOfShapeListOfShape from TopTools,
    Edge from TopoDS, Shape from TopoDS

is

    Create returns EdgeConnect from ShapeFix;

    Add (me : in out; aFirst : Edge from TopoDS; aSecond : Edge from TopoDS);
    ---Purpose : Adds information on connectivity between start vertex
    --           of second edge and end vertex of first edge,
    --           taking edges orientation into account

    Add (me : in out; aShape : Shape from TopoDS);
    ---Purpose : Adds connectivity information for the whole shape.
    --           Note: edges in wires must be well ordered
    --           Note: flag Closed should be set for closed wires

    Build (me : in out);
    ---Purpose : Builds shared vertices, updates their positions and tolerances

    Clear (me : in out);
    ---Purpose : Clears internal data structure

fields

    myVertices : DataMapOfShapeShape from TopTools;       -- Map of pairs (vertex, shared)
    myLists    : DataMapOfShapeListOfShape from TopTools; -- Map of pairs (shared, list of vertices/edges)

end EdgeConnect;
